magic
tech sky130A
timestamp 1701310363
<< locali >>
rect 24 131 41 162
rect 133 -27 150 29
rect -15 -44 189 -27
rect -141 -333 -124 -270
rect 298 -332 315 -271
rect -32 -548 -15 -537
rect 189 -547 206 -536
use sky130_fd_pr__nfet_01v8_8BU2MY  sky130_fd_pr__nfet_01v8_8BU2MY_0
timestamp 1701309485
transform 1 0 252 0 1 -434
box -69 -113 69 113
use sky130_fd_pr__nfet_01v8_8BU2MY  sky130_fd_pr__nfet_01v8_8BU2MY_1
timestamp 1701309485
transform 1 0 -78 0 1 -435
box -69 -113 69 113
use sky130_fd_pr__pfet_01v8_ES6STC  sky130_fd_pr__pfet_01v8_ES6STC_0
timestamp 1701309268
transform 1 0 87 0 1 81
box -87 -81 87 81
use sky130_fd_pr__pfet_01v8_S43UTC  sky130_fd_pr__pfet_01v8_S43UTC_0
timestamp 1701309268
transform 1 0 252 0 1 -69
box -87 -231 87 231
use sky130_fd_pr__pfet_01v8_S43UTC  sky130_fd_pr__pfet_01v8_S43UTC_1
timestamp 1701309268
transform 1 0 -78 0 1 -69
box -87 -231 87 231
<< end >>

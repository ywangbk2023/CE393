* NGSPICE file created from SARLOGIC_layout.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
**devattr s=8216,420 d=4582,216
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
**devattr s=3016,162 d=5408,312
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
**devattr s=4582,216 d=8216,420
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
**devattr s=5408,312 d=3016,162
.ends

.subckt sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 a_788_47# a_942_21# a_648_21# VNB sky130_fd_pr__nfet_01v8 ad=0.139 pd=1.42 as=0.0864 ps=0.91 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X1 VPWR RESET_B a_942_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.16 as=0.166 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6156,267
X2 VGND a_1429_21# a_1364_47# VNB sky130_fd_pr__nfet_01v8 ad=0.078 pd=0.843 as=0.0711 ps=0.802 w=0.42 l=0.15
**devattr s=2640,149 d=2352,140
X3 VPWR a_942_21# a_1663_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.53 as=0.0882 ps=1.05 w=0.84 l=0.15
**devattr s=3528,210 d=8736,440
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.16 as=0.166 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.086 ps=0.763 w=0.42 l=0.15
**devattr s=4368,272 d=2646,147
X6 VPWR a_1429_21# a_1341_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.086 pd=0.763 as=0.0924 ps=0.86 w=0.42 l=0.15
**devattr s=3696,172 d=3276,162
X7 a_474_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.0609 ps=0.688 w=0.36 l=0.15
**devattr s=2640,149 d=2736,148
X8 a_1545_47# a_942_21# a_1429_21# VNB sky130_fd_pr__nfet_01v8 ad=0.153 pd=1.49 as=0.0864 ps=0.91 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X9 VPWR a_1429_21# a_2136_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.131 pd=1.16 as=0.166 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=5960,265
X10 a_582_47# a_193_47# a_474_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0619 pd=0.692 as=0.0684 ps=0.74 w=0.36 l=0.15
**devattr s=2736,148 d=2682,150
X11 a_1429_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.78 as=0.086 ps=0.763 w=0.42 l=0.15
**devattr s=3276,162 d=4914,234
X12 a_648_21# a_474_413# a_788_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.139 ps=1.42 w=0.64 l=0.15
**devattr s=4040,198 d=3456,182
X13 a_1341_413# a_193_47# a_1255_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3696,172
X14 a_1663_329# a_1255_47# a_1429_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.164 ps=1.56 w=0.84 l=0.15
**devattr s=4914,234 d=3528,210
X15 a_1160_47# a_648_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.24 as=0.119 ps=1.28 w=0.64 l=0.15
**devattr s=6656,360 d=3740,193
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.078 ps=0.843 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X17 a_1255_47# a_27_47# a_1113_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.116 ps=0.94 w=0.42 l=0.15
**devattr s=6972,282 d=2268,138
X18 Q a_2136_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.205 ps=1.82 w=1 l=0.15
**devattr s=5960,265 d=10400,504
X19 a_648_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.098 pd=0.82 as=0.086 ps=0.763 w=0.42 l=0.15
**devattr s=3192,160 d=5880,246
X20 a_788_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.934 as=0.078 ps=0.843 w=0.42 l=0.15
**devattr s=3360,164 d=4040,198
X21 Q_N a_1429_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.205 ps=1.82 w=1 l=0.15
**devattr s=6156,267 d=10400,504
X22 VGND RESET_B a_942_21# VNB sky130_fd_pr__nfet_01v8 ad=0.078 pd=0.843 as=0.109 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X23 Q a_2136_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.121 ps=1.3 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X24 VPWR a_942_21# a_892_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.53 as=0.113 ps=1.11 w=0.84 l=0.15
**devattr s=4536,222 d=8988,275
X25 a_558_413# a_27_47# a_474_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3780,174
X26 VGND a_648_21# a_582_47# VNB sky130_fd_pr__nfet_01v8 ad=0.078 pd=0.843 as=0.0722 ps=0.808 w=0.42 l=0.15
**devattr s=2682,150 d=3360,164
X27 a_892_329# a_474_413# a_648_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.196 ps=1.64 w=0.84 l=0.15
**devattr s=5880,246 d=4536,222
X28 VGND a_1429_21# a_2136_47# VNB sky130_fd_pr__nfet_01v8 ad=0.078 pd=0.843 as=0.109 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=3880,195
X29 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.131 ps=1.16 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X30 a_474_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
**devattr s=2646,147 d=2268,138
X31 a_1364_47# a_27_47# a_1255_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.688 as=0.0711 ps=0.755 w=0.36 l=0.15
**devattr s=2844,151 d=2640,149
X32 a_1255_47# a_193_47# a_1160_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0673 ps=0.695 w=0.36 l=0.15
**devattr s=3740,193 d=2844,151
X33 Q_N a_1429_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.121 ps=1.3 w=0.65 l=0.15
**devattr s=3880,195 d=6760,364
X34 a_1545_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.978 as=0.078 ps=0.843 w=0.42 l=0.15
**devattr s=2352,140 d=4796,216
X35 VPWR a_648_21# a_558_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.086 pd=0.763 as=0.0945 ps=0.87 w=0.42 l=0.15
**devattr s=3780,174 d=3192,160
X36 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.802 as=0.078 ps=0.843 w=0.42 l=0.15
**devattr s=4368,272 d=2640,149
X37 a_1113_329# a_648_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.232 pd=1.88 as=0.172 ps=1.53 w=0.84 l=0.15
**devattr s=8988,275 d=6972,282
X38 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.078 pd=0.843 as=0.109 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X39 a_1429_21# a_1255_47# a_1545_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.153 ps=1.49 w=0.64 l=0.15
**devattr s=4796,216 d=3456,182
.ends

.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N a_1847_47#
+ a_27_47#
X0 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.211 ps=1.99 w=1 l=0.15
**devattr s=8528,334 d=11200,512
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0618 pd=0.692 as=0.0711 ps=0.755 w=0.36 l=0.15
**devattr s=2844,151 d=2676,150
X2 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.151 ps=1.18 w=0.42 l=0.15
**devattr s=5604,220 d=1764,126
X3 VPWR a_1283_21# a_1847_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.28 as=0.166 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=6160,267
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0719 ps=0.709 w=0.36 l=0.15
**devattr s=3996,197 d=2844,151
X5 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
**devattr s=2562,145 d=4368,272
X6 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.1 as=0.0724 ps=0.765 w=0.42 l=0.15
**devattr s=2898,153 d=4620,194
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.98 as=0.0441 ps=0.63 w=0.42 l=0.15
**devattr s=1764,126 d=5384,230
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.28 as=0.166 ps=1.8 w=0.64 l=0.15
**devattr s=6656,360 d=3456,182
X9 Q_N a_1847_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.163 ps=1.52 w=0.65 l=0.15
**devattr s=4010,197 d=6760,364
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.0888 ps=0.838 w=0.42 l=0.15
**devattr s=4368,272 d=2604,146
X11 VGND a_1283_21# a_1847_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.98 as=0.109 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=4010,197
X12 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.128 pd=1.26 as=0.16 ps=1.49 w=0.64 l=0.15
**devattr s=5384,230 d=3996,197
X13 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.163 ps=1.52 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.105 ps=0.98 w=0.42 l=0.15
**devattr s=2268,138 d=4368,272
X15 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0861 ps=0.79 w=0.42 l=0.15
**devattr s=5166,237 d=2352,140
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.0609 ps=0.688 w=0.36 l=0.15
**devattr s=2640,149 d=2376,138
X17 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.105 ps=0.98 w=0.42 l=0.15
**devattr s=4998,203 d=2562,145
X18 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
**devattr s=2604,146 d=2898,153
X19 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.802 as=0.105 ps=0.98 w=0.42 l=0.15
**devattr s=8820,378 d=2640,149
X20 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0888 pd=0.838 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=3276,162
X21 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0888 pd=0.838 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=8528,334
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
**devattr s=2352,140 d=2268,138
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.135 ps=1.28 w=0.64 l=0.15
**devattr s=3456,182 d=6656,360
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0888 ps=0.838 w=0.42 l=0.15
**devattr s=3276,162 d=2268,138
X25 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0888 pd=0.838 as=0.113 ps=1.1 w=0.42 l=0.15
**devattr s=4620,194 d=2814,151
X26 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.129 pd=1.02 as=0.0594 ps=0.69 w=0.36 l=0.15
**devattr s=2376,138 d=5604,220
X27 Q_N a_1847_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.211 ps=1.99 w=1 l=0.15
**devattr s=6160,267 d=10400,504
X28 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.98 as=0.072 ps=0.808 w=0.42 l=0.15
**devattr s=2676,150 d=4998,203
X29 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.1 as=0.0888 ps=0.838 w=0.42 l=0.15
**devattr s=2814,151 d=4368,272
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.105 pd=0.98 as=0.109 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2268,138
X31 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.58 as=0.178 ps=1.68 w=0.84 l=0.15
**devattr s=8736,440 d=5166,237
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=6760,364
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
.ends

.subckt SARLOGIC_layout dout6 dout5 dout4 doutb4 dout1 dout3 dout2
Xsky130_fd_sc_hd__buf_1_4 sky130_fd_sc_hd__buf_1_4/A sky130_fd_sc_hd__inv_1_0/VGND
+ VSUBS sky130_fd_sc_hd__inv_1_0/VPB sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__buf_1_4/X
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__dfbbp_1_0 sky130_fd_sc_hd__dfbbp_1_5/Q sky130_fd_sc_hd__buf_1_2/X
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__dfrbp_1_6/Q_N sky130_fd_sc_hd__dfrbp_1_8/VGND
+ VSUBS sky130_fd_sc_hd__dfbbp_1_7/VPB sky130_fd_sc_hd__dfbbp_1_7/VPWR dout1 sky130_fd_sc_hd__dfbbp_1_0/Q_N
+ sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_1 dout5 sky130_fd_sc_hd__buf_1_2/X sky130_fd_sc_hd__buf_1_3/X
+ sky130_fd_sc_hd__dfrbp_1_2/Q_N sky130_fd_sc_hd__inv_1_0/VGND VSUBS sky130_fd_sc_hd__buf_1_2/VPB
+ sky130_fd_sc_hd__buf_1_2/VPWR dout6 sky130_fd_sc_hd__dfbbp_1_1/Q_N sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_2 dout4 sky130_fd_sc_hd__buf_1_2/X sky130_fd_sc_hd__buf_1_3/X
+ sky130_fd_sc_hd__dfrbp_1_1/Q_N sky130_fd_sc_hd__inv_1_0/VGND VSUBS sky130_fd_sc_hd__buf_1_2/VPB
+ sky130_fd_sc_hd__buf_1_2/VPWR dout5 sky130_fd_sc_hd__dfbbp_1_2/Q_N sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_3 sky130_fd_sc_hd__dfbbp_1_3/CLK sky130_fd_sc_hd__buf_1_2/X
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__dfrbp_1_3/Q_N sky130_fd_sc_hd__inv_1_0/VGND
+ VSUBS sky130_fd_sc_hd__buf_1_2/VPB sky130_fd_sc_hd__buf_1_2/VPWR dout4 sky130_fd_sc_hd__dfbbp_1_3/Q_N
+ sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_4 dout6 sky130_fd_sc_hd__buf_1_2/X sky130_fd_sc_hd__buf_1_3/X
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__inv_1_0/VGND VSUBS sky130_fd_sc_hd__buf_1_2/VPB
+ sky130_fd_sc_hd__buf_1_2/VPWR sky130_fd_sc_hd__dfbbp_1_4/Q sky130_fd_sc_hd__dfbbp_1_4/Q_N
+ sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_6 dout1 sky130_fd_sc_hd__buf_1_2/X sky130_fd_sc_hd__buf_1_3/X
+ sky130_fd_sc_hd__dfrbp_1_7/Q_N sky130_fd_sc_hd__dfrbp_1_8/VGND VSUBS sky130_fd_sc_hd__dfbbp_1_7/VPB
+ sky130_fd_sc_hd__dfbbp_1_7/VPWR sky130_fd_sc_hd__dfbbp_1_6/Q sky130_fd_sc_hd__dfbbp_1_6/Q_N
+ sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_5 sky130_fd_sc_hd__dfrbp_1_8/Q sky130_fd_sc_hd__buf_1_2/X
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__dfrbp_1_5/Q_N sky130_fd_sc_hd__dfrbp_1_8/VGND
+ VSUBS sky130_fd_sc_hd__dfbbp_1_7/VPB sky130_fd_sc_hd__dfbbp_1_7/VPWR sky130_fd_sc_hd__dfbbp_1_5/Q
+ sky130_fd_sc_hd__dfbbp_1_5/Q_N sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_7 dout2 sky130_fd_sc_hd__buf_1_2/X sky130_fd_sc_hd__buf_1_3/X
+ sky130_fd_sc_hd__dfrbp_1_4/Q_N sky130_fd_sc_hd__dfrbp_1_8/VGND VSUBS sky130_fd_sc_hd__dfbbp_1_7/VPB
+ sky130_fd_sc_hd__dfbbp_1_7/VPWR dout3 sky130_fd_sc_hd__dfbbp_1_7/Q_N sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfrbp_1_0 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__buf_1_0/X
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__inv_1_0/VGND VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__dfrbp_1_2/D sky130_fd_sc_hd__buf_1_3/X
+ sky130_fd_sc_hd__dfrbp_1_0/a_1847_47# sky130_fd_sc_hd__buf_1_0/X sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_1 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__dfrbp_1_2/Q
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__inv_1_0/VGND VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__dfrbp_1_3/D sky130_fd_sc_hd__dfrbp_1_1/Q_N
+ sky130_fd_sc_hd__dfrbp_1_1/a_1847_47# sky130_fd_sc_hd__dfrbp_1_1/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_2 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__dfrbp_1_2/D
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__inv_1_0/VGND VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__dfrbp_1_2/Q sky130_fd_sc_hd__dfrbp_1_2/Q_N
+ sky130_fd_sc_hd__dfrbp_1_2/a_1847_47# sky130_fd_sc_hd__dfrbp_1_2/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_3 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__dfrbp_1_3/D
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__inv_1_0/VGND VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__dfrbp_1_4/D sky130_fd_sc_hd__dfrbp_1_3/Q_N
+ sky130_fd_sc_hd__dfrbp_1_3/a_1847_47# sky130_fd_sc_hd__dfrbp_1_3/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_4 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__dfrbp_1_4/D
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__dfrbp_1_8/VGND VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__dfrbp_1_7/D sky130_fd_sc_hd__dfrbp_1_4/Q_N
+ sky130_fd_sc_hd__dfrbp_1_4/a_1847_47# sky130_fd_sc_hd__dfrbp_1_4/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_5 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__dfrbp_1_6/Q
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__dfrbp_1_8/VGND VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__dfrbp_1_5/Q sky130_fd_sc_hd__dfrbp_1_5/Q_N
+ sky130_fd_sc_hd__dfrbp_1_8/D sky130_fd_sc_hd__dfrbp_1_5/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_6 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__dfrbp_1_7/Q
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__dfrbp_1_8/VGND VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__dfrbp_1_6/Q sky130_fd_sc_hd__dfrbp_1_6/Q_N
+ sky130_fd_sc_hd__dfrbp_1_6/a_1847_47# sky130_fd_sc_hd__dfrbp_1_6/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_7 sky130_fd_sc_hd__inv_1_0/Y sky130_fd_sc_hd__dfrbp_1_7/D
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__dfrbp_1_8/VGND VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__dfrbp_1_7/Q sky130_fd_sc_hd__dfrbp_1_7/Q_N
+ sky130_fd_sc_hd__dfrbp_1_7/a_1847_47# sky130_fd_sc_hd__dfrbp_1_7/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__buf_1_0 sky130_fd_sc_hd__buf_1_0/A sky130_fd_sc_hd__inv_1_0/VGND
+ VSUBS sky130_fd_sc_hd__inv_1_0/VPB sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__buf_1_0/X
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__dfrbp_1_8 sky130_fd_sc_hd__dfrbp_1_8/CLK sky130_fd_sc_hd__dfrbp_1_8/D
+ sky130_fd_sc_hd__buf_1_3/X sky130_fd_sc_hd__dfrbp_1_8/VGND VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__dfrbp_1_8/Q sky130_fd_sc_hd__dfrbp_1_8/Q_N
+ sky130_fd_sc_hd__dfrbp_1_8/a_1847_47# sky130_fd_sc_hd__dfrbp_1_8/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/A sky130_fd_sc_hd__inv_1_0/VGND
+ VSUBS sky130_fd_sc_hd__inv_1_0/VPB sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__inv_1_0/Y
+ sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__buf_1_1 sky130_fd_sc_hd__buf_1_1/A sky130_fd_sc_hd__inv_1_0/VGND
+ VSUBS sky130_fd_sc_hd__inv_1_0/VPB sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__inv_1_0/A
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_2 sky130_fd_sc_hd__buf_1_2/A sky130_fd_sc_hd__inv_1_0/VGND
+ VSUBS sky130_fd_sc_hd__buf_1_2/VPB sky130_fd_sc_hd__buf_1_2/VPWR sky130_fd_sc_hd__buf_1_2/X
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_3 sky130_fd_sc_hd__buf_1_4/X sky130_fd_sc_hd__inv_1_0/VGND
+ VSUBS sky130_fd_sc_hd__inv_1_0/VPB sky130_fd_sc_hd__inv_1_0/VPWR sky130_fd_sc_hd__buf_1_3/X
+ sky130_fd_sc_hd__buf_1
.ends


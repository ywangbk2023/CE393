magic
tech sky130A
magscale 1 2
timestamp 1701908128
<< metal3 >>
rect -29634 12492 -23262 12520
rect -29634 6468 -23346 12492
rect -23282 6468 -23262 12492
rect -29634 6440 -23262 6468
rect -23022 12492 -16650 12520
rect -23022 6468 -16734 12492
rect -16670 6468 -16650 12492
rect -23022 6440 -16650 6468
rect -16410 12492 -10038 12520
rect -16410 6468 -10122 12492
rect -10058 6468 -10038 12492
rect -16410 6440 -10038 6468
rect -9798 12492 -3426 12520
rect -9798 6468 -3510 12492
rect -3446 6468 -3426 12492
rect -9798 6440 -3426 6468
rect -3186 12492 3186 12520
rect -3186 6468 3102 12492
rect 3166 6468 3186 12492
rect -3186 6440 3186 6468
rect 3426 12492 9798 12520
rect 3426 6468 9714 12492
rect 9778 6468 9798 12492
rect 3426 6440 9798 6468
rect 10038 12492 16410 12520
rect 10038 6468 16326 12492
rect 16390 6468 16410 12492
rect 10038 6440 16410 6468
rect 16650 12492 23022 12520
rect 16650 6468 22938 12492
rect 23002 6468 23022 12492
rect 16650 6440 23022 6468
rect 23262 12492 29634 12520
rect 23262 6468 29550 12492
rect 29614 6468 29634 12492
rect 23262 6440 29634 6468
rect -29634 6172 -23262 6200
rect -29634 148 -23346 6172
rect -23282 148 -23262 6172
rect -29634 120 -23262 148
rect -23022 6172 -16650 6200
rect -23022 148 -16734 6172
rect -16670 148 -16650 6172
rect -23022 120 -16650 148
rect -16410 6172 -10038 6200
rect -16410 148 -10122 6172
rect -10058 148 -10038 6172
rect -16410 120 -10038 148
rect -9798 6172 -3426 6200
rect -9798 148 -3510 6172
rect -3446 148 -3426 6172
rect -9798 120 -3426 148
rect -3186 6172 3186 6200
rect -3186 148 3102 6172
rect 3166 148 3186 6172
rect -3186 120 3186 148
rect 3426 6172 9798 6200
rect 3426 148 9714 6172
rect 9778 148 9798 6172
rect 3426 120 9798 148
rect 10038 6172 16410 6200
rect 10038 148 16326 6172
rect 16390 148 16410 6172
rect 10038 120 16410 148
rect 16650 6172 23022 6200
rect 16650 148 22938 6172
rect 23002 148 23022 6172
rect 16650 120 23022 148
rect 23262 6172 29634 6200
rect 23262 148 29550 6172
rect 29614 148 29634 6172
rect 23262 120 29634 148
rect -29634 -148 -23262 -120
rect -29634 -6172 -23346 -148
rect -23282 -6172 -23262 -148
rect -29634 -6200 -23262 -6172
rect -23022 -148 -16650 -120
rect -23022 -6172 -16734 -148
rect -16670 -6172 -16650 -148
rect -23022 -6200 -16650 -6172
rect -16410 -148 -10038 -120
rect -16410 -6172 -10122 -148
rect -10058 -6172 -10038 -148
rect -16410 -6200 -10038 -6172
rect -9798 -148 -3426 -120
rect -9798 -6172 -3510 -148
rect -3446 -6172 -3426 -148
rect -9798 -6200 -3426 -6172
rect -3186 -148 3186 -120
rect -3186 -6172 3102 -148
rect 3166 -6172 3186 -148
rect -3186 -6200 3186 -6172
rect 3426 -148 9798 -120
rect 3426 -6172 9714 -148
rect 9778 -6172 9798 -148
rect 3426 -6200 9798 -6172
rect 10038 -148 16410 -120
rect 10038 -6172 16326 -148
rect 16390 -6172 16410 -148
rect 10038 -6200 16410 -6172
rect 16650 -148 23022 -120
rect 16650 -6172 22938 -148
rect 23002 -6172 23022 -148
rect 16650 -6200 23022 -6172
rect 23262 -148 29634 -120
rect 23262 -6172 29550 -148
rect 29614 -6172 29634 -148
rect 23262 -6200 29634 -6172
rect -29634 -6468 -23262 -6440
rect -29634 -12492 -23346 -6468
rect -23282 -12492 -23262 -6468
rect -29634 -12520 -23262 -12492
rect -23022 -6468 -16650 -6440
rect -23022 -12492 -16734 -6468
rect -16670 -12492 -16650 -6468
rect -23022 -12520 -16650 -12492
rect -16410 -6468 -10038 -6440
rect -16410 -12492 -10122 -6468
rect -10058 -12492 -10038 -6468
rect -16410 -12520 -10038 -12492
rect -9798 -6468 -3426 -6440
rect -9798 -12492 -3510 -6468
rect -3446 -12492 -3426 -6468
rect -9798 -12520 -3426 -12492
rect -3186 -6468 3186 -6440
rect -3186 -12492 3102 -6468
rect 3166 -12492 3186 -6468
rect -3186 -12520 3186 -12492
rect 3426 -6468 9798 -6440
rect 3426 -12492 9714 -6468
rect 9778 -12492 9798 -6468
rect 3426 -12520 9798 -12492
rect 10038 -6468 16410 -6440
rect 10038 -12492 16326 -6468
rect 16390 -12492 16410 -6468
rect 10038 -12520 16410 -12492
rect 16650 -6468 23022 -6440
rect 16650 -12492 22938 -6468
rect 23002 -12492 23022 -6468
rect 16650 -12520 23022 -12492
rect 23262 -6468 29634 -6440
rect 23262 -12492 29550 -6468
rect 29614 -12492 29634 -6468
rect 23262 -12520 29634 -12492
<< via3 >>
rect -23346 6468 -23282 12492
rect -16734 6468 -16670 12492
rect -10122 6468 -10058 12492
rect -3510 6468 -3446 12492
rect 3102 6468 3166 12492
rect 9714 6468 9778 12492
rect 16326 6468 16390 12492
rect 22938 6468 23002 12492
rect 29550 6468 29614 12492
rect -23346 148 -23282 6172
rect -16734 148 -16670 6172
rect -10122 148 -10058 6172
rect -3510 148 -3446 6172
rect 3102 148 3166 6172
rect 9714 148 9778 6172
rect 16326 148 16390 6172
rect 22938 148 23002 6172
rect 29550 148 29614 6172
rect -23346 -6172 -23282 -148
rect -16734 -6172 -16670 -148
rect -10122 -6172 -10058 -148
rect -3510 -6172 -3446 -148
rect 3102 -6172 3166 -148
rect 9714 -6172 9778 -148
rect 16326 -6172 16390 -148
rect 22938 -6172 23002 -148
rect 29550 -6172 29614 -148
rect -23346 -12492 -23282 -6468
rect -16734 -12492 -16670 -6468
rect -10122 -12492 -10058 -6468
rect -3510 -12492 -3446 -6468
rect 3102 -12492 3166 -6468
rect 9714 -12492 9778 -6468
rect 16326 -12492 16390 -6468
rect 22938 -12492 23002 -6468
rect 29550 -12492 29614 -6468
<< mimcap >>
rect -29594 12440 -23594 12480
rect -29594 6520 -29554 12440
rect -23634 6520 -23594 12440
rect -29594 6480 -23594 6520
rect -22982 12440 -16982 12480
rect -22982 6520 -22942 12440
rect -17022 6520 -16982 12440
rect -22982 6480 -16982 6520
rect -16370 12440 -10370 12480
rect -16370 6520 -16330 12440
rect -10410 6520 -10370 12440
rect -16370 6480 -10370 6520
rect -9758 12440 -3758 12480
rect -9758 6520 -9718 12440
rect -3798 6520 -3758 12440
rect -9758 6480 -3758 6520
rect -3146 12440 2854 12480
rect -3146 6520 -3106 12440
rect 2814 6520 2854 12440
rect -3146 6480 2854 6520
rect 3466 12440 9466 12480
rect 3466 6520 3506 12440
rect 9426 6520 9466 12440
rect 3466 6480 9466 6520
rect 10078 12440 16078 12480
rect 10078 6520 10118 12440
rect 16038 6520 16078 12440
rect 10078 6480 16078 6520
rect 16690 12440 22690 12480
rect 16690 6520 16730 12440
rect 22650 6520 22690 12440
rect 16690 6480 22690 6520
rect 23302 12440 29302 12480
rect 23302 6520 23342 12440
rect 29262 6520 29302 12440
rect 23302 6480 29302 6520
rect -29594 6120 -23594 6160
rect -29594 200 -29554 6120
rect -23634 200 -23594 6120
rect -29594 160 -23594 200
rect -22982 6120 -16982 6160
rect -22982 200 -22942 6120
rect -17022 200 -16982 6120
rect -22982 160 -16982 200
rect -16370 6120 -10370 6160
rect -16370 200 -16330 6120
rect -10410 200 -10370 6120
rect -16370 160 -10370 200
rect -9758 6120 -3758 6160
rect -9758 200 -9718 6120
rect -3798 200 -3758 6120
rect -9758 160 -3758 200
rect -3146 6120 2854 6160
rect -3146 200 -3106 6120
rect 2814 200 2854 6120
rect -3146 160 2854 200
rect 3466 6120 9466 6160
rect 3466 200 3506 6120
rect 9426 200 9466 6120
rect 3466 160 9466 200
rect 10078 6120 16078 6160
rect 10078 200 10118 6120
rect 16038 200 16078 6120
rect 10078 160 16078 200
rect 16690 6120 22690 6160
rect 16690 200 16730 6120
rect 22650 200 22690 6120
rect 16690 160 22690 200
rect 23302 6120 29302 6160
rect 23302 200 23342 6120
rect 29262 200 29302 6120
rect 23302 160 29302 200
rect -29594 -200 -23594 -160
rect -29594 -6120 -29554 -200
rect -23634 -6120 -23594 -200
rect -29594 -6160 -23594 -6120
rect -22982 -200 -16982 -160
rect -22982 -6120 -22942 -200
rect -17022 -6120 -16982 -200
rect -22982 -6160 -16982 -6120
rect -16370 -200 -10370 -160
rect -16370 -6120 -16330 -200
rect -10410 -6120 -10370 -200
rect -16370 -6160 -10370 -6120
rect -9758 -200 -3758 -160
rect -9758 -6120 -9718 -200
rect -3798 -6120 -3758 -200
rect -9758 -6160 -3758 -6120
rect -3146 -200 2854 -160
rect -3146 -6120 -3106 -200
rect 2814 -6120 2854 -200
rect -3146 -6160 2854 -6120
rect 3466 -200 9466 -160
rect 3466 -6120 3506 -200
rect 9426 -6120 9466 -200
rect 3466 -6160 9466 -6120
rect 10078 -200 16078 -160
rect 10078 -6120 10118 -200
rect 16038 -6120 16078 -200
rect 10078 -6160 16078 -6120
rect 16690 -200 22690 -160
rect 16690 -6120 16730 -200
rect 22650 -6120 22690 -200
rect 16690 -6160 22690 -6120
rect 23302 -200 29302 -160
rect 23302 -6120 23342 -200
rect 29262 -6120 29302 -200
rect 23302 -6160 29302 -6120
rect -29594 -6520 -23594 -6480
rect -29594 -12440 -29554 -6520
rect -23634 -12440 -23594 -6520
rect -29594 -12480 -23594 -12440
rect -22982 -6520 -16982 -6480
rect -22982 -12440 -22942 -6520
rect -17022 -12440 -16982 -6520
rect -22982 -12480 -16982 -12440
rect -16370 -6520 -10370 -6480
rect -16370 -12440 -16330 -6520
rect -10410 -12440 -10370 -6520
rect -16370 -12480 -10370 -12440
rect -9758 -6520 -3758 -6480
rect -9758 -12440 -9718 -6520
rect -3798 -12440 -3758 -6520
rect -9758 -12480 -3758 -12440
rect -3146 -6520 2854 -6480
rect -3146 -12440 -3106 -6520
rect 2814 -12440 2854 -6520
rect -3146 -12480 2854 -12440
rect 3466 -6520 9466 -6480
rect 3466 -12440 3506 -6520
rect 9426 -12440 9466 -6520
rect 3466 -12480 9466 -12440
rect 10078 -6520 16078 -6480
rect 10078 -12440 10118 -6520
rect 16038 -12440 16078 -6520
rect 10078 -12480 16078 -12440
rect 16690 -6520 22690 -6480
rect 16690 -12440 16730 -6520
rect 22650 -12440 22690 -6520
rect 16690 -12480 22690 -12440
rect 23302 -6520 29302 -6480
rect 23302 -12440 23342 -6520
rect 29262 -12440 29302 -6520
rect 23302 -12480 29302 -12440
<< mimcapcontact >>
rect -29554 6520 -23634 12440
rect -22942 6520 -17022 12440
rect -16330 6520 -10410 12440
rect -9718 6520 -3798 12440
rect -3106 6520 2814 12440
rect 3506 6520 9426 12440
rect 10118 6520 16038 12440
rect 16730 6520 22650 12440
rect 23342 6520 29262 12440
rect -29554 200 -23634 6120
rect -22942 200 -17022 6120
rect -16330 200 -10410 6120
rect -9718 200 -3798 6120
rect -3106 200 2814 6120
rect 3506 200 9426 6120
rect 10118 200 16038 6120
rect 16730 200 22650 6120
rect 23342 200 29262 6120
rect -29554 -6120 -23634 -200
rect -22942 -6120 -17022 -200
rect -16330 -6120 -10410 -200
rect -9718 -6120 -3798 -200
rect -3106 -6120 2814 -200
rect 3506 -6120 9426 -200
rect 10118 -6120 16038 -200
rect 16730 -6120 22650 -200
rect 23342 -6120 29262 -200
rect -29554 -12440 -23634 -6520
rect -22942 -12440 -17022 -6520
rect -16330 -12440 -10410 -6520
rect -9718 -12440 -3798 -6520
rect -3106 -12440 2814 -6520
rect 3506 -12440 9426 -6520
rect 10118 -12440 16038 -6520
rect 16730 -12440 22650 -6520
rect 23342 -12440 29262 -6520
<< metal4 >>
rect -26646 12441 -26542 12640
rect -23366 12492 -23262 12640
rect -29555 12440 -23633 12441
rect -29555 6520 -29554 12440
rect -23634 6520 -23633 12440
rect -29555 6519 -23633 6520
rect -26646 6121 -26542 6519
rect -23366 6468 -23346 12492
rect -23282 6468 -23262 12492
rect -20034 12441 -19930 12640
rect -16754 12492 -16650 12640
rect -22943 12440 -17021 12441
rect -22943 6520 -22942 12440
rect -17022 6520 -17021 12440
rect -22943 6519 -17021 6520
rect -23366 6172 -23262 6468
rect -29555 6120 -23633 6121
rect -29555 200 -29554 6120
rect -23634 200 -23633 6120
rect -29555 199 -23633 200
rect -26646 -199 -26542 199
rect -23366 148 -23346 6172
rect -23282 148 -23262 6172
rect -20034 6121 -19930 6519
rect -16754 6468 -16734 12492
rect -16670 6468 -16650 12492
rect -13422 12441 -13318 12640
rect -10142 12492 -10038 12640
rect -16331 12440 -10409 12441
rect -16331 6520 -16330 12440
rect -10410 6520 -10409 12440
rect -16331 6519 -10409 6520
rect -16754 6172 -16650 6468
rect -22943 6120 -17021 6121
rect -22943 200 -22942 6120
rect -17022 200 -17021 6120
rect -22943 199 -17021 200
rect -23366 -148 -23262 148
rect -29555 -200 -23633 -199
rect -29555 -6120 -29554 -200
rect -23634 -6120 -23633 -200
rect -29555 -6121 -23633 -6120
rect -26646 -6519 -26542 -6121
rect -23366 -6172 -23346 -148
rect -23282 -6172 -23262 -148
rect -20034 -199 -19930 199
rect -16754 148 -16734 6172
rect -16670 148 -16650 6172
rect -13422 6121 -13318 6519
rect -10142 6468 -10122 12492
rect -10058 6468 -10038 12492
rect -6810 12441 -6706 12640
rect -3530 12492 -3426 12640
rect -9719 12440 -3797 12441
rect -9719 6520 -9718 12440
rect -3798 6520 -3797 12440
rect -9719 6519 -3797 6520
rect -10142 6172 -10038 6468
rect -16331 6120 -10409 6121
rect -16331 200 -16330 6120
rect -10410 200 -10409 6120
rect -16331 199 -10409 200
rect -16754 -148 -16650 148
rect -22943 -200 -17021 -199
rect -22943 -6120 -22942 -200
rect -17022 -6120 -17021 -200
rect -22943 -6121 -17021 -6120
rect -23366 -6468 -23262 -6172
rect -29555 -6520 -23633 -6519
rect -29555 -12440 -29554 -6520
rect -23634 -12440 -23633 -6520
rect -29555 -12441 -23633 -12440
rect -26646 -12640 -26542 -12441
rect -23366 -12492 -23346 -6468
rect -23282 -12492 -23262 -6468
rect -20034 -6519 -19930 -6121
rect -16754 -6172 -16734 -148
rect -16670 -6172 -16650 -148
rect -13422 -199 -13318 199
rect -10142 148 -10122 6172
rect -10058 148 -10038 6172
rect -6810 6121 -6706 6519
rect -3530 6468 -3510 12492
rect -3446 6468 -3426 12492
rect -198 12441 -94 12640
rect 3082 12492 3186 12640
rect -3107 12440 2815 12441
rect -3107 6520 -3106 12440
rect 2814 6520 2815 12440
rect -3107 6519 2815 6520
rect -3530 6172 -3426 6468
rect -9719 6120 -3797 6121
rect -9719 200 -9718 6120
rect -3798 200 -3797 6120
rect -9719 199 -3797 200
rect -10142 -148 -10038 148
rect -16331 -200 -10409 -199
rect -16331 -6120 -16330 -200
rect -10410 -6120 -10409 -200
rect -16331 -6121 -10409 -6120
rect -16754 -6468 -16650 -6172
rect -22943 -6520 -17021 -6519
rect -22943 -12440 -22942 -6520
rect -17022 -12440 -17021 -6520
rect -22943 -12441 -17021 -12440
rect -23366 -12640 -23262 -12492
rect -20034 -12640 -19930 -12441
rect -16754 -12492 -16734 -6468
rect -16670 -12492 -16650 -6468
rect -13422 -6519 -13318 -6121
rect -10142 -6172 -10122 -148
rect -10058 -6172 -10038 -148
rect -6810 -199 -6706 199
rect -3530 148 -3510 6172
rect -3446 148 -3426 6172
rect -198 6121 -94 6519
rect 3082 6468 3102 12492
rect 3166 6468 3186 12492
rect 6414 12441 6518 12640
rect 9694 12492 9798 12640
rect 3505 12440 9427 12441
rect 3505 6520 3506 12440
rect 9426 6520 9427 12440
rect 3505 6519 9427 6520
rect 3082 6172 3186 6468
rect -3107 6120 2815 6121
rect -3107 200 -3106 6120
rect 2814 200 2815 6120
rect -3107 199 2815 200
rect -3530 -148 -3426 148
rect -9719 -200 -3797 -199
rect -9719 -6120 -9718 -200
rect -3798 -6120 -3797 -200
rect -9719 -6121 -3797 -6120
rect -10142 -6468 -10038 -6172
rect -16331 -6520 -10409 -6519
rect -16331 -12440 -16330 -6520
rect -10410 -12440 -10409 -6520
rect -16331 -12441 -10409 -12440
rect -16754 -12640 -16650 -12492
rect -13422 -12640 -13318 -12441
rect -10142 -12492 -10122 -6468
rect -10058 -12492 -10038 -6468
rect -6810 -6519 -6706 -6121
rect -3530 -6172 -3510 -148
rect -3446 -6172 -3426 -148
rect -198 -199 -94 199
rect 3082 148 3102 6172
rect 3166 148 3186 6172
rect 6414 6121 6518 6519
rect 9694 6468 9714 12492
rect 9778 6468 9798 12492
rect 13026 12441 13130 12640
rect 16306 12492 16410 12640
rect 10117 12440 16039 12441
rect 10117 6520 10118 12440
rect 16038 6520 16039 12440
rect 10117 6519 16039 6520
rect 9694 6172 9798 6468
rect 3505 6120 9427 6121
rect 3505 200 3506 6120
rect 9426 200 9427 6120
rect 3505 199 9427 200
rect 3082 -148 3186 148
rect -3107 -200 2815 -199
rect -3107 -6120 -3106 -200
rect 2814 -6120 2815 -200
rect -3107 -6121 2815 -6120
rect -3530 -6468 -3426 -6172
rect -9719 -6520 -3797 -6519
rect -9719 -12440 -9718 -6520
rect -3798 -12440 -3797 -6520
rect -9719 -12441 -3797 -12440
rect -10142 -12640 -10038 -12492
rect -6810 -12640 -6706 -12441
rect -3530 -12492 -3510 -6468
rect -3446 -12492 -3426 -6468
rect -198 -6519 -94 -6121
rect 3082 -6172 3102 -148
rect 3166 -6172 3186 -148
rect 6414 -199 6518 199
rect 9694 148 9714 6172
rect 9778 148 9798 6172
rect 13026 6121 13130 6519
rect 16306 6468 16326 12492
rect 16390 6468 16410 12492
rect 19638 12441 19742 12640
rect 22918 12492 23022 12640
rect 16729 12440 22651 12441
rect 16729 6520 16730 12440
rect 22650 6520 22651 12440
rect 16729 6519 22651 6520
rect 16306 6172 16410 6468
rect 10117 6120 16039 6121
rect 10117 200 10118 6120
rect 16038 200 16039 6120
rect 10117 199 16039 200
rect 9694 -148 9798 148
rect 3505 -200 9427 -199
rect 3505 -6120 3506 -200
rect 9426 -6120 9427 -200
rect 3505 -6121 9427 -6120
rect 3082 -6468 3186 -6172
rect -3107 -6520 2815 -6519
rect -3107 -12440 -3106 -6520
rect 2814 -12440 2815 -6520
rect -3107 -12441 2815 -12440
rect -3530 -12640 -3426 -12492
rect -198 -12640 -94 -12441
rect 3082 -12492 3102 -6468
rect 3166 -12492 3186 -6468
rect 6414 -6519 6518 -6121
rect 9694 -6172 9714 -148
rect 9778 -6172 9798 -148
rect 13026 -199 13130 199
rect 16306 148 16326 6172
rect 16390 148 16410 6172
rect 19638 6121 19742 6519
rect 22918 6468 22938 12492
rect 23002 6468 23022 12492
rect 26250 12441 26354 12640
rect 29530 12492 29634 12640
rect 23341 12440 29263 12441
rect 23341 6520 23342 12440
rect 29262 6520 29263 12440
rect 23341 6519 29263 6520
rect 22918 6172 23022 6468
rect 16729 6120 22651 6121
rect 16729 200 16730 6120
rect 22650 200 22651 6120
rect 16729 199 22651 200
rect 16306 -148 16410 148
rect 10117 -200 16039 -199
rect 10117 -6120 10118 -200
rect 16038 -6120 16039 -200
rect 10117 -6121 16039 -6120
rect 9694 -6468 9798 -6172
rect 3505 -6520 9427 -6519
rect 3505 -12440 3506 -6520
rect 9426 -12440 9427 -6520
rect 3505 -12441 9427 -12440
rect 3082 -12640 3186 -12492
rect 6414 -12640 6518 -12441
rect 9694 -12492 9714 -6468
rect 9778 -12492 9798 -6468
rect 13026 -6519 13130 -6121
rect 16306 -6172 16326 -148
rect 16390 -6172 16410 -148
rect 19638 -199 19742 199
rect 22918 148 22938 6172
rect 23002 148 23022 6172
rect 26250 6121 26354 6519
rect 29530 6468 29550 12492
rect 29614 6468 29634 12492
rect 29530 6172 29634 6468
rect 23341 6120 29263 6121
rect 23341 200 23342 6120
rect 29262 200 29263 6120
rect 23341 199 29263 200
rect 22918 -148 23022 148
rect 16729 -200 22651 -199
rect 16729 -6120 16730 -200
rect 22650 -6120 22651 -200
rect 16729 -6121 22651 -6120
rect 16306 -6468 16410 -6172
rect 10117 -6520 16039 -6519
rect 10117 -12440 10118 -6520
rect 16038 -12440 16039 -6520
rect 10117 -12441 16039 -12440
rect 9694 -12640 9798 -12492
rect 13026 -12640 13130 -12441
rect 16306 -12492 16326 -6468
rect 16390 -12492 16410 -6468
rect 19638 -6519 19742 -6121
rect 22918 -6172 22938 -148
rect 23002 -6172 23022 -148
rect 26250 -199 26354 199
rect 29530 148 29550 6172
rect 29614 148 29634 6172
rect 29530 -148 29634 148
rect 23341 -200 29263 -199
rect 23341 -6120 23342 -200
rect 29262 -6120 29263 -200
rect 23341 -6121 29263 -6120
rect 22918 -6468 23022 -6172
rect 16729 -6520 22651 -6519
rect 16729 -12440 16730 -6520
rect 22650 -12440 22651 -6520
rect 16729 -12441 22651 -12440
rect 16306 -12640 16410 -12492
rect 19638 -12640 19742 -12441
rect 22918 -12492 22938 -6468
rect 23002 -12492 23022 -6468
rect 26250 -6519 26354 -6121
rect 29530 -6172 29550 -148
rect 29614 -6172 29634 -148
rect 29530 -6468 29634 -6172
rect 23341 -6520 29263 -6519
rect 23341 -12440 23342 -6520
rect 29262 -12440 29263 -6520
rect 23341 -12441 29263 -12440
rect 22918 -12640 23022 -12492
rect 26250 -12640 26354 -12441
rect 29530 -12492 29550 -6468
rect 29614 -12492 29634 -6468
rect 29530 -12640 29634 -12492
<< properties >>
string FIXED_BBOX 23262 6440 29342 12520
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 9 ny 4 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

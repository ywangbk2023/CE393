magic
tech sky130A
magscale 1 2
timestamp 1702102630
<< error_s >>
rect 577 1079 590 1103
rect 611 1045 624 1069
rect 966 1035 1001 1069
rect 967 1016 1001 1035
rect 775 967 837 973
rect 775 933 787 967
rect 775 927 837 933
rect 276 813 317 819
rect 575 599 584 797
rect 775 623 837 629
rect 577 535 590 569
rect 611 501 624 603
rect 775 589 787 623
rect 775 583 837 589
rect 986 487 1001 1016
rect 1020 982 1055 1016
rect 1020 487 1054 982
rect 1184 914 1246 920
rect 1184 880 1196 914
rect 1184 874 1246 880
rect 1184 570 1246 576
rect 1184 536 1196 570
rect 1184 530 1246 536
rect 1020 453 1035 487
rect 1395 434 1410 1016
rect 1429 434 1463 1070
rect 1593 1019 1655 1025
rect 1593 985 1605 1019
rect 1593 979 1655 985
rect 1785 910 1819 964
rect 1593 517 1655 523
rect 1593 483 1605 517
rect 1593 477 1655 483
rect 1429 400 1444 434
rect 1804 381 1819 910
rect 1838 876 1873 910
rect 2193 876 2228 910
rect 1838 381 1872 876
rect 2194 857 2228 876
rect 2002 808 2064 814
rect 2002 774 2014 808
rect 2002 768 2064 774
rect 2002 464 2064 470
rect 2002 430 2014 464
rect 2002 424 2064 430
rect 1838 347 1853 381
rect 2213 328 2228 857
rect 2247 823 2282 857
rect 2247 328 2281 823
rect 2411 755 2473 761
rect 2411 721 2423 755
rect 2411 715 2473 721
rect 2411 411 2473 417
rect 2411 377 2423 411
rect 2411 371 2473 377
rect 2247 294 2262 328
rect 2622 275 2637 857
rect 2656 275 2690 911
rect 2820 860 2882 866
rect 2820 826 2832 860
rect 2820 820 2882 826
rect 3012 673 3046 691
rect 3012 637 3082 673
rect 3029 603 3100 637
rect 3380 603 3415 637
rect 2820 358 2882 364
rect 2820 324 2832 358
rect 2820 318 2882 324
rect 2656 241 2671 275
rect 3029 222 3099 603
rect 3381 584 3415 603
rect 3211 535 3269 541
rect 3211 501 3223 535
rect 3211 495 3269 501
rect 3211 305 3269 311
rect 3211 271 3223 305
rect 3211 265 3269 271
rect 3029 186 3082 222
rect 3400 169 3415 584
rect 3434 550 3469 584
rect 3749 550 3784 584
rect 3434 169 3468 550
rect 3750 531 3784 550
rect 3580 482 3638 488
rect 3580 448 3592 482
rect 3580 442 3638 448
rect 3580 252 3638 258
rect 3580 218 3592 252
rect 3580 212 3638 218
rect 3434 135 3449 169
rect 3769 116 3784 531
rect 3803 497 3838 531
rect 4118 497 4153 531
rect 3803 116 3837 497
rect 4119 478 4153 497
rect 3949 429 4007 435
rect 3949 395 3961 429
rect 3949 389 4007 395
rect 3949 199 4007 205
rect 3949 165 3961 199
rect 3949 159 4007 165
rect 3803 82 3818 116
rect 4138 63 4153 478
rect 4172 444 4207 478
rect 4487 444 4522 478
rect 4172 63 4206 444
rect 4488 425 4522 444
rect 4318 376 4376 382
rect 4318 342 4330 376
rect 4318 336 4376 342
rect 4318 146 4376 152
rect 4318 112 4330 146
rect 4318 106 4376 112
rect 4172 29 4187 63
rect 4507 10 4522 425
rect 4541 391 4576 425
rect 4541 10 4575 391
rect 4687 323 4745 329
rect 4687 289 4699 323
rect 4687 283 4745 289
rect 4687 93 4745 99
rect 4687 59 4699 93
rect 4687 53 4745 59
rect 4541 -24 4556 10
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
rect 0 -1200 200 -1000
rect 0 -1600 200 -1400
rect 0 -2000 200 -1800
use sky130_fd_sc_hd__buf_1  x1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697562905
transform 1 0 0 0 1 600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  x2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697562905
transform 1 0 314 0 1 552
box -38 -48 314 592
use sky130_fd_pr__pfet_01v8_NFJWV9  XM1
timestamp 1702102630
transform 1 0 806 0 1 778
box -231 -327 231 327
use sky130_fd_pr__pfet_01v8_NFJWV9  XM2
timestamp 1702102630
transform 1 0 1215 0 1 725
box -231 -327 231 327
use sky130_fd_pr__pfet_01v8_NFFSV9  XM3
timestamp 1702102630
transform 1 0 1624 0 1 751
box -231 -406 231 406
use sky130_fd_pr__pfet_01v8_NFJWV9  XM4
timestamp 1702102630
transform 1 0 2033 0 1 619
box -231 -327 231 327
use sky130_fd_pr__pfet_01v8_NFJWV9  XM5
timestamp 1702102630
transform 1 0 2442 0 1 566
box -231 -327 231 327
use sky130_fd_pr__pfet_01v8_NFFSV9  XM6
timestamp 1702102630
transform 1 0 2851 0 1 592
box -231 -406 231 406
use sky130_fd_pr__nfet_01v8_HNLS78  XM7
timestamp 1702102630
transform 1 0 3240 0 1 403
box -211 -270 211 270
use sky130_fd_pr__nfet_01v8_HNLS78  XM8
timestamp 1702102630
transform 1 0 3609 0 1 350
box -211 -270 211 270
use sky130_fd_pr__nfet_01v8_HNLS78  XM9
timestamp 1702102630
transform 1 0 3978 0 1 297
box -211 -270 211 270
use sky130_fd_pr__nfet_01v8_HNLS78  XM10
timestamp 1702102630
transform 1 0 4347 0 1 244
box -211 -270 211 270
use sky130_fd_pr__nfet_01v8_HNLS78  XM11
timestamp 1702102630
transform 1 0 4716 0 1 191
box -211 -270 211 270
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VSS
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VDD
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Vref
port 2 nsew
flabel metal1 0 -1200 200 -1000 0 FreeSans 256 0 0 0 Vmac
port 3 nsew
flabel metal1 0 -1600 200 -1400 0 FreeSans 256 0 0 0 Clk
port 4 nsew
flabel metal1 0 -2000 200 -1800 0 FreeSans 256 0 0 0 Updown
port 5 nsew
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1701405958
<< error_p >>
rect -29 399 29 405
rect -29 365 -17 399
rect -29 359 29 365
rect -29 71 29 77
rect -29 37 -17 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect -29 -77 29 -71
rect -29 -365 29 -359
rect -29 -399 -17 -365
rect -29 -405 29 -399
<< nwell >>
rect -211 -537 211 537
<< pmos >>
rect -15 118 15 318
rect -15 -318 15 -118
<< pdiff >>
rect -73 306 -15 318
rect -73 130 -61 306
rect -27 130 -15 306
rect -73 118 -15 130
rect 15 306 73 318
rect 15 130 27 306
rect 61 130 73 306
rect 15 118 73 130
rect -73 -130 -15 -118
rect -73 -306 -61 -130
rect -27 -306 -15 -130
rect -73 -318 -15 -306
rect 15 -130 73 -118
rect 15 -306 27 -130
rect 61 -306 73 -130
rect 15 -318 73 -306
<< pdiffc >>
rect -61 130 -27 306
rect 27 130 61 306
rect -61 -306 -27 -130
rect 27 -306 61 -130
<< nsubdiff >>
rect -175 467 -79 501
rect 79 467 175 501
rect -175 405 -141 467
rect 141 405 175 467
rect -175 -467 -141 -405
rect 141 -467 175 -405
rect -175 -501 -79 -467
rect 79 -501 175 -467
<< nsubdiffcont >>
rect -79 467 79 501
rect -175 -405 -141 405
rect 141 -405 175 405
rect -79 -501 79 -467
<< poly >>
rect -33 399 33 415
rect -33 365 -17 399
rect 17 365 33 399
rect -33 349 33 365
rect -15 318 15 349
rect -15 87 15 118
rect -33 71 33 87
rect -33 37 -17 71
rect 17 37 33 71
rect -33 21 33 37
rect -33 -37 33 -21
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -33 -87 33 -71
rect -15 -118 15 -87
rect -15 -349 15 -318
rect -33 -365 33 -349
rect -33 -399 -17 -365
rect 17 -399 33 -365
rect -33 -415 33 -399
<< polycont >>
rect -17 365 17 399
rect -17 37 17 71
rect -17 -71 17 -37
rect -17 -399 17 -365
<< locali >>
rect -175 467 -79 501
rect 79 467 175 501
rect -175 405 -141 467
rect 141 405 175 467
rect -33 365 -17 399
rect 17 365 33 399
rect -61 306 -27 322
rect -61 114 -27 130
rect 27 306 61 322
rect 27 114 61 130
rect -33 37 -17 71
rect 17 37 33 71
rect -33 -71 -17 -37
rect 17 -71 33 -37
rect -61 -130 -27 -114
rect -61 -322 -27 -306
rect 27 -130 61 -114
rect 27 -322 61 -306
rect -33 -399 -17 -365
rect 17 -399 33 -365
rect -175 -467 -141 -405
rect 141 -467 175 -405
rect -175 -501 -79 -467
rect 79 -501 175 -467
<< viali >>
rect -17 365 17 399
rect -61 130 -27 306
rect 27 130 61 306
rect -17 37 17 71
rect -17 -71 17 -37
rect -61 -306 -27 -130
rect 27 -306 61 -130
rect -17 -399 17 -365
<< metal1 >>
rect -29 399 29 405
rect -29 365 -17 399
rect 17 365 29 399
rect -29 359 29 365
rect -67 306 -21 318
rect -67 130 -61 306
rect -27 130 -21 306
rect -67 118 -21 130
rect 21 306 67 318
rect 21 130 27 306
rect 61 130 67 306
rect 21 118 67 130
rect -29 71 29 77
rect -29 37 -17 71
rect 17 37 29 71
rect -29 31 29 37
rect -29 -37 29 -31
rect -29 -71 -17 -37
rect 17 -71 29 -37
rect -29 -77 29 -71
rect -67 -130 -21 -118
rect -67 -306 -61 -130
rect -27 -306 -21 -130
rect -67 -318 -21 -306
rect 21 -130 67 -118
rect 21 -306 27 -130
rect 61 -306 67 -130
rect 21 -318 67 -306
rect -29 -365 29 -359
rect -29 -399 -17 -365
rect 17 -399 29 -365
rect -29 -405 29 -399
<< properties >>
string FIXED_BBOX -158 -484 158 484
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 2 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1701909930
<< metal3 >>
rect -19710 18806 -13340 18834
rect -19710 12784 -13424 18806
rect -13360 12784 -13340 18806
rect -19710 12756 -13340 12784
rect -13100 18806 -6730 18834
rect -13100 12784 -6814 18806
rect -6750 12784 -6730 18806
rect -13100 12756 -6730 12784
rect -6490 18806 -120 18834
rect -6490 12784 -204 18806
rect -140 12784 -120 18806
rect -6490 12756 -120 12784
rect 120 18806 6490 18834
rect 120 12784 6406 18806
rect 6470 12784 6490 18806
rect 120 12756 6490 12784
rect 6730 18806 13100 18834
rect 6730 12784 13016 18806
rect 13080 12784 13100 18806
rect 6730 12756 13100 12784
rect 13340 18806 19710 18834
rect 13340 12784 19626 18806
rect 19690 12784 19710 18806
rect 13340 12756 19710 12784
rect -19710 12488 -13340 12516
rect -19710 6466 -13424 12488
rect -13360 6466 -13340 12488
rect -19710 6438 -13340 6466
rect -13100 12488 -6730 12516
rect -13100 6466 -6814 12488
rect -6750 6466 -6730 12488
rect -13100 6438 -6730 6466
rect -6490 12488 -120 12516
rect -6490 6466 -204 12488
rect -140 6466 -120 12488
rect -6490 6438 -120 6466
rect 120 12488 6490 12516
rect 120 6466 6406 12488
rect 6470 6466 6490 12488
rect 120 6438 6490 6466
rect 6730 12488 13100 12516
rect 6730 6466 13016 12488
rect 13080 6466 13100 12488
rect 6730 6438 13100 6466
rect 13340 12488 19710 12516
rect 13340 6466 19626 12488
rect 19690 6466 19710 12488
rect 13340 6438 19710 6466
rect -19710 6170 -13340 6198
rect -19710 148 -13424 6170
rect -13360 148 -13340 6170
rect -19710 120 -13340 148
rect -13100 6170 -6730 6198
rect -13100 148 -6814 6170
rect -6750 148 -6730 6170
rect -13100 120 -6730 148
rect -6490 6170 -120 6198
rect -6490 148 -204 6170
rect -140 148 -120 6170
rect -6490 120 -120 148
rect 120 6170 6490 6198
rect 120 148 6406 6170
rect 6470 148 6490 6170
rect 120 120 6490 148
rect 6730 6170 13100 6198
rect 6730 148 13016 6170
rect 13080 148 13100 6170
rect 6730 120 13100 148
rect 13340 6170 19710 6198
rect 13340 148 19626 6170
rect 19690 148 19710 6170
rect 13340 120 19710 148
rect -19710 -148 -13340 -120
rect -19710 -6170 -13424 -148
rect -13360 -6170 -13340 -148
rect -19710 -6198 -13340 -6170
rect -13100 -148 -6730 -120
rect -13100 -6170 -6814 -148
rect -6750 -6170 -6730 -148
rect -13100 -6198 -6730 -6170
rect -6490 -148 -120 -120
rect -6490 -6170 -204 -148
rect -140 -6170 -120 -148
rect -6490 -6198 -120 -6170
rect 120 -148 6490 -120
rect 120 -6170 6406 -148
rect 6470 -6170 6490 -148
rect 120 -6198 6490 -6170
rect 6730 -148 13100 -120
rect 6730 -6170 13016 -148
rect 13080 -6170 13100 -148
rect 6730 -6198 13100 -6170
rect 13340 -148 19710 -120
rect 13340 -6170 19626 -148
rect 19690 -6170 19710 -148
rect 13340 -6198 19710 -6170
rect -19710 -6466 -13340 -6438
rect -19710 -12488 -13424 -6466
rect -13360 -12488 -13340 -6466
rect -19710 -12516 -13340 -12488
rect -13100 -6466 -6730 -6438
rect -13100 -12488 -6814 -6466
rect -6750 -12488 -6730 -6466
rect -13100 -12516 -6730 -12488
rect -6490 -6466 -120 -6438
rect -6490 -12488 -204 -6466
rect -140 -12488 -120 -6466
rect -6490 -12516 -120 -12488
rect 120 -6466 6490 -6438
rect 120 -12488 6406 -6466
rect 6470 -12488 6490 -6466
rect 120 -12516 6490 -12488
rect 6730 -6466 13100 -6438
rect 6730 -12488 13016 -6466
rect 13080 -12488 13100 -6466
rect 6730 -12516 13100 -12488
rect 13340 -6466 19710 -6438
rect 13340 -12488 19626 -6466
rect 19690 -12488 19710 -6466
rect 13340 -12516 19710 -12488
rect -19710 -12784 -13340 -12756
rect -19710 -18806 -13424 -12784
rect -13360 -18806 -13340 -12784
rect -19710 -18834 -13340 -18806
rect -13100 -12784 -6730 -12756
rect -13100 -18806 -6814 -12784
rect -6750 -18806 -6730 -12784
rect -13100 -18834 -6730 -18806
rect -6490 -12784 -120 -12756
rect -6490 -18806 -204 -12784
rect -140 -18806 -120 -12784
rect -6490 -18834 -120 -18806
rect 120 -12784 6490 -12756
rect 120 -18806 6406 -12784
rect 6470 -18806 6490 -12784
rect 120 -18834 6490 -18806
rect 6730 -12784 13100 -12756
rect 6730 -18806 13016 -12784
rect 13080 -18806 13100 -12784
rect 6730 -18834 13100 -18806
rect 13340 -12784 19710 -12756
rect 13340 -18806 19626 -12784
rect 19690 -18806 19710 -12784
rect 13340 -18834 19710 -18806
<< via3 >>
rect -13424 12784 -13360 18806
rect -6814 12784 -6750 18806
rect -204 12784 -140 18806
rect 6406 12784 6470 18806
rect 13016 12784 13080 18806
rect 19626 12784 19690 18806
rect -13424 6466 -13360 12488
rect -6814 6466 -6750 12488
rect -204 6466 -140 12488
rect 6406 6466 6470 12488
rect 13016 6466 13080 12488
rect 19626 6466 19690 12488
rect -13424 148 -13360 6170
rect -6814 148 -6750 6170
rect -204 148 -140 6170
rect 6406 148 6470 6170
rect 13016 148 13080 6170
rect 19626 148 19690 6170
rect -13424 -6170 -13360 -148
rect -6814 -6170 -6750 -148
rect -204 -6170 -140 -148
rect 6406 -6170 6470 -148
rect 13016 -6170 13080 -148
rect 19626 -6170 19690 -148
rect -13424 -12488 -13360 -6466
rect -6814 -12488 -6750 -6466
rect -204 -12488 -140 -6466
rect 6406 -12488 6470 -6466
rect 13016 -12488 13080 -6466
rect 19626 -12488 19690 -6466
rect -13424 -18806 -13360 -12784
rect -6814 -18806 -6750 -12784
rect -204 -18806 -140 -12784
rect 6406 -18806 6470 -12784
rect 13016 -18806 13080 -12784
rect 19626 -18806 19690 -12784
<< mimcap >>
rect -19670 18754 -13672 18794
rect -19670 12836 -19630 18754
rect -13712 12836 -13672 18754
rect -19670 12796 -13672 12836
rect -13060 18754 -7062 18794
rect -13060 12836 -13020 18754
rect -7102 12836 -7062 18754
rect -13060 12796 -7062 12836
rect -6450 18754 -452 18794
rect -6450 12836 -6410 18754
rect -492 12836 -452 18754
rect -6450 12796 -452 12836
rect 160 18754 6158 18794
rect 160 12836 200 18754
rect 6118 12836 6158 18754
rect 160 12796 6158 12836
rect 6770 18754 12768 18794
rect 6770 12836 6810 18754
rect 12728 12836 12768 18754
rect 6770 12796 12768 12836
rect 13380 18754 19378 18794
rect 13380 12836 13420 18754
rect 19338 12836 19378 18754
rect 13380 12796 19378 12836
rect -19670 12436 -13672 12476
rect -19670 6518 -19630 12436
rect -13712 6518 -13672 12436
rect -19670 6478 -13672 6518
rect -13060 12436 -7062 12476
rect -13060 6518 -13020 12436
rect -7102 6518 -7062 12436
rect -13060 6478 -7062 6518
rect -6450 12436 -452 12476
rect -6450 6518 -6410 12436
rect -492 6518 -452 12436
rect -6450 6478 -452 6518
rect 160 12436 6158 12476
rect 160 6518 200 12436
rect 6118 6518 6158 12436
rect 160 6478 6158 6518
rect 6770 12436 12768 12476
rect 6770 6518 6810 12436
rect 12728 6518 12768 12436
rect 6770 6478 12768 6518
rect 13380 12436 19378 12476
rect 13380 6518 13420 12436
rect 19338 6518 19378 12436
rect 13380 6478 19378 6518
rect -19670 6118 -13672 6158
rect -19670 200 -19630 6118
rect -13712 200 -13672 6118
rect -19670 160 -13672 200
rect -13060 6118 -7062 6158
rect -13060 200 -13020 6118
rect -7102 200 -7062 6118
rect -13060 160 -7062 200
rect -6450 6118 -452 6158
rect -6450 200 -6410 6118
rect -492 200 -452 6118
rect -6450 160 -452 200
rect 160 6118 6158 6158
rect 160 200 200 6118
rect 6118 200 6158 6118
rect 160 160 6158 200
rect 6770 6118 12768 6158
rect 6770 200 6810 6118
rect 12728 200 12768 6118
rect 6770 160 12768 200
rect 13380 6118 19378 6158
rect 13380 200 13420 6118
rect 19338 200 19378 6118
rect 13380 160 19378 200
rect -19670 -200 -13672 -160
rect -19670 -6118 -19630 -200
rect -13712 -6118 -13672 -200
rect -19670 -6158 -13672 -6118
rect -13060 -200 -7062 -160
rect -13060 -6118 -13020 -200
rect -7102 -6118 -7062 -200
rect -13060 -6158 -7062 -6118
rect -6450 -200 -452 -160
rect -6450 -6118 -6410 -200
rect -492 -6118 -452 -200
rect -6450 -6158 -452 -6118
rect 160 -200 6158 -160
rect 160 -6118 200 -200
rect 6118 -6118 6158 -200
rect 160 -6158 6158 -6118
rect 6770 -200 12768 -160
rect 6770 -6118 6810 -200
rect 12728 -6118 12768 -200
rect 6770 -6158 12768 -6118
rect 13380 -200 19378 -160
rect 13380 -6118 13420 -200
rect 19338 -6118 19378 -200
rect 13380 -6158 19378 -6118
rect -19670 -6518 -13672 -6478
rect -19670 -12436 -19630 -6518
rect -13712 -12436 -13672 -6518
rect -19670 -12476 -13672 -12436
rect -13060 -6518 -7062 -6478
rect -13060 -12436 -13020 -6518
rect -7102 -12436 -7062 -6518
rect -13060 -12476 -7062 -12436
rect -6450 -6518 -452 -6478
rect -6450 -12436 -6410 -6518
rect -492 -12436 -452 -6518
rect -6450 -12476 -452 -12436
rect 160 -6518 6158 -6478
rect 160 -12436 200 -6518
rect 6118 -12436 6158 -6518
rect 160 -12476 6158 -12436
rect 6770 -6518 12768 -6478
rect 6770 -12436 6810 -6518
rect 12728 -12436 12768 -6518
rect 6770 -12476 12768 -12436
rect 13380 -6518 19378 -6478
rect 13380 -12436 13420 -6518
rect 19338 -12436 19378 -6518
rect 13380 -12476 19378 -12436
rect -19670 -12836 -13672 -12796
rect -19670 -18754 -19630 -12836
rect -13712 -18754 -13672 -12836
rect -19670 -18794 -13672 -18754
rect -13060 -12836 -7062 -12796
rect -13060 -18754 -13020 -12836
rect -7102 -18754 -7062 -12836
rect -13060 -18794 -7062 -18754
rect -6450 -12836 -452 -12796
rect -6450 -18754 -6410 -12836
rect -492 -18754 -452 -12836
rect -6450 -18794 -452 -18754
rect 160 -12836 6158 -12796
rect 160 -18754 200 -12836
rect 6118 -18754 6158 -12836
rect 160 -18794 6158 -18754
rect 6770 -12836 12768 -12796
rect 6770 -18754 6810 -12836
rect 12728 -18754 12768 -12836
rect 6770 -18794 12768 -18754
rect 13380 -12836 19378 -12796
rect 13380 -18754 13420 -12836
rect 19338 -18754 19378 -12836
rect 13380 -18794 19378 -18754
<< mimcapcontact >>
rect -19630 12836 -13712 18754
rect -13020 12836 -7102 18754
rect -6410 12836 -492 18754
rect 200 12836 6118 18754
rect 6810 12836 12728 18754
rect 13420 12836 19338 18754
rect -19630 6518 -13712 12436
rect -13020 6518 -7102 12436
rect -6410 6518 -492 12436
rect 200 6518 6118 12436
rect 6810 6518 12728 12436
rect 13420 6518 19338 12436
rect -19630 200 -13712 6118
rect -13020 200 -7102 6118
rect -6410 200 -492 6118
rect 200 200 6118 6118
rect 6810 200 12728 6118
rect 13420 200 19338 6118
rect -19630 -6118 -13712 -200
rect -13020 -6118 -7102 -200
rect -6410 -6118 -492 -200
rect 200 -6118 6118 -200
rect 6810 -6118 12728 -200
rect 13420 -6118 19338 -200
rect -19630 -12436 -13712 -6518
rect -13020 -12436 -7102 -6518
rect -6410 -12436 -492 -6518
rect 200 -12436 6118 -6518
rect 6810 -12436 12728 -6518
rect 13420 -12436 19338 -6518
rect -19630 -18754 -13712 -12836
rect -13020 -18754 -7102 -12836
rect -6410 -18754 -492 -12836
rect 200 -18754 6118 -12836
rect 6810 -18754 12728 -12836
rect 13420 -18754 19338 -12836
<< metal4 >>
rect -16723 18755 -16619 18954
rect -13444 18806 -13340 18954
rect -19631 18754 -13711 18755
rect -19631 12836 -19630 18754
rect -13712 12836 -13711 18754
rect -19631 12835 -13711 12836
rect -16723 12437 -16619 12835
rect -13444 12784 -13424 18806
rect -13360 12784 -13340 18806
rect -10113 18755 -10009 18954
rect -6834 18806 -6730 18954
rect -13021 18754 -7101 18755
rect -13021 12836 -13020 18754
rect -7102 12836 -7101 18754
rect -13021 12835 -7101 12836
rect -13444 12488 -13340 12784
rect -19631 12436 -13711 12437
rect -19631 6518 -19630 12436
rect -13712 6518 -13711 12436
rect -19631 6517 -13711 6518
rect -16723 6119 -16619 6517
rect -13444 6466 -13424 12488
rect -13360 6466 -13340 12488
rect -10113 12437 -10009 12835
rect -6834 12784 -6814 18806
rect -6750 12784 -6730 18806
rect -3503 18755 -3399 18954
rect -224 18806 -120 18954
rect -6411 18754 -491 18755
rect -6411 12836 -6410 18754
rect -492 12836 -491 18754
rect -6411 12835 -491 12836
rect -6834 12488 -6730 12784
rect -13021 12436 -7101 12437
rect -13021 6518 -13020 12436
rect -7102 6518 -7101 12436
rect -13021 6517 -7101 6518
rect -13444 6170 -13340 6466
rect -19631 6118 -13711 6119
rect -19631 200 -19630 6118
rect -13712 200 -13711 6118
rect -19631 199 -13711 200
rect -16723 -199 -16619 199
rect -13444 148 -13424 6170
rect -13360 148 -13340 6170
rect -10113 6119 -10009 6517
rect -6834 6466 -6814 12488
rect -6750 6466 -6730 12488
rect -3503 12437 -3399 12835
rect -224 12784 -204 18806
rect -140 12784 -120 18806
rect 3107 18755 3211 18954
rect 6386 18806 6490 18954
rect 199 18754 6119 18755
rect 199 12836 200 18754
rect 6118 12836 6119 18754
rect 199 12835 6119 12836
rect -224 12488 -120 12784
rect -6411 12436 -491 12437
rect -6411 6518 -6410 12436
rect -492 6518 -491 12436
rect -6411 6517 -491 6518
rect -6834 6170 -6730 6466
rect -13021 6118 -7101 6119
rect -13021 200 -13020 6118
rect -7102 200 -7101 6118
rect -13021 199 -7101 200
rect -13444 -148 -13340 148
rect -19631 -200 -13711 -199
rect -19631 -6118 -19630 -200
rect -13712 -6118 -13711 -200
rect -19631 -6119 -13711 -6118
rect -16723 -6517 -16619 -6119
rect -13444 -6170 -13424 -148
rect -13360 -6170 -13340 -148
rect -10113 -199 -10009 199
rect -6834 148 -6814 6170
rect -6750 148 -6730 6170
rect -3503 6119 -3399 6517
rect -224 6466 -204 12488
rect -140 6466 -120 12488
rect 3107 12437 3211 12835
rect 6386 12784 6406 18806
rect 6470 12784 6490 18806
rect 9717 18755 9821 18954
rect 12996 18806 13100 18954
rect 6809 18754 12729 18755
rect 6809 12836 6810 18754
rect 12728 12836 12729 18754
rect 6809 12835 12729 12836
rect 6386 12488 6490 12784
rect 199 12436 6119 12437
rect 199 6518 200 12436
rect 6118 6518 6119 12436
rect 199 6517 6119 6518
rect -224 6170 -120 6466
rect -6411 6118 -491 6119
rect -6411 200 -6410 6118
rect -492 200 -491 6118
rect -6411 199 -491 200
rect -6834 -148 -6730 148
rect -13021 -200 -7101 -199
rect -13021 -6118 -13020 -200
rect -7102 -6118 -7101 -200
rect -13021 -6119 -7101 -6118
rect -13444 -6466 -13340 -6170
rect -19631 -6518 -13711 -6517
rect -19631 -12436 -19630 -6518
rect -13712 -12436 -13711 -6518
rect -19631 -12437 -13711 -12436
rect -16723 -12835 -16619 -12437
rect -13444 -12488 -13424 -6466
rect -13360 -12488 -13340 -6466
rect -10113 -6517 -10009 -6119
rect -6834 -6170 -6814 -148
rect -6750 -6170 -6730 -148
rect -3503 -199 -3399 199
rect -224 148 -204 6170
rect -140 148 -120 6170
rect 3107 6119 3211 6517
rect 6386 6466 6406 12488
rect 6470 6466 6490 12488
rect 9717 12437 9821 12835
rect 12996 12784 13016 18806
rect 13080 12784 13100 18806
rect 16327 18755 16431 18954
rect 19606 18806 19710 18954
rect 13419 18754 19339 18755
rect 13419 12836 13420 18754
rect 19338 12836 19339 18754
rect 13419 12835 19339 12836
rect 12996 12488 13100 12784
rect 6809 12436 12729 12437
rect 6809 6518 6810 12436
rect 12728 6518 12729 12436
rect 6809 6517 12729 6518
rect 6386 6170 6490 6466
rect 199 6118 6119 6119
rect 199 200 200 6118
rect 6118 200 6119 6118
rect 199 199 6119 200
rect -224 -148 -120 148
rect -6411 -200 -491 -199
rect -6411 -6118 -6410 -200
rect -492 -6118 -491 -200
rect -6411 -6119 -491 -6118
rect -6834 -6466 -6730 -6170
rect -13021 -6518 -7101 -6517
rect -13021 -12436 -13020 -6518
rect -7102 -12436 -7101 -6518
rect -13021 -12437 -7101 -12436
rect -13444 -12784 -13340 -12488
rect -19631 -12836 -13711 -12835
rect -19631 -18754 -19630 -12836
rect -13712 -18754 -13711 -12836
rect -19631 -18755 -13711 -18754
rect -16723 -18954 -16619 -18755
rect -13444 -18806 -13424 -12784
rect -13360 -18806 -13340 -12784
rect -10113 -12835 -10009 -12437
rect -6834 -12488 -6814 -6466
rect -6750 -12488 -6730 -6466
rect -3503 -6517 -3399 -6119
rect -224 -6170 -204 -148
rect -140 -6170 -120 -148
rect 3107 -199 3211 199
rect 6386 148 6406 6170
rect 6470 148 6490 6170
rect 9717 6119 9821 6517
rect 12996 6466 13016 12488
rect 13080 6466 13100 12488
rect 16327 12437 16431 12835
rect 19606 12784 19626 18806
rect 19690 12784 19710 18806
rect 19606 12488 19710 12784
rect 13419 12436 19339 12437
rect 13419 6518 13420 12436
rect 19338 6518 19339 12436
rect 13419 6517 19339 6518
rect 12996 6170 13100 6466
rect 6809 6118 12729 6119
rect 6809 200 6810 6118
rect 12728 200 12729 6118
rect 6809 199 12729 200
rect 6386 -148 6490 148
rect 199 -200 6119 -199
rect 199 -6118 200 -200
rect 6118 -6118 6119 -200
rect 199 -6119 6119 -6118
rect -224 -6466 -120 -6170
rect -6411 -6518 -491 -6517
rect -6411 -12436 -6410 -6518
rect -492 -12436 -491 -6518
rect -6411 -12437 -491 -12436
rect -6834 -12784 -6730 -12488
rect -13021 -12836 -7101 -12835
rect -13021 -18754 -13020 -12836
rect -7102 -18754 -7101 -12836
rect -13021 -18755 -7101 -18754
rect -13444 -18954 -13340 -18806
rect -10113 -18954 -10009 -18755
rect -6834 -18806 -6814 -12784
rect -6750 -18806 -6730 -12784
rect -3503 -12835 -3399 -12437
rect -224 -12488 -204 -6466
rect -140 -12488 -120 -6466
rect 3107 -6517 3211 -6119
rect 6386 -6170 6406 -148
rect 6470 -6170 6490 -148
rect 9717 -199 9821 199
rect 12996 148 13016 6170
rect 13080 148 13100 6170
rect 16327 6119 16431 6517
rect 19606 6466 19626 12488
rect 19690 6466 19710 12488
rect 19606 6170 19710 6466
rect 13419 6118 19339 6119
rect 13419 200 13420 6118
rect 19338 200 19339 6118
rect 13419 199 19339 200
rect 12996 -148 13100 148
rect 6809 -200 12729 -199
rect 6809 -6118 6810 -200
rect 12728 -6118 12729 -200
rect 6809 -6119 12729 -6118
rect 6386 -6466 6490 -6170
rect 199 -6518 6119 -6517
rect 199 -12436 200 -6518
rect 6118 -12436 6119 -6518
rect 199 -12437 6119 -12436
rect -224 -12784 -120 -12488
rect -6411 -12836 -491 -12835
rect -6411 -18754 -6410 -12836
rect -492 -18754 -491 -12836
rect -6411 -18755 -491 -18754
rect -6834 -18954 -6730 -18806
rect -3503 -18954 -3399 -18755
rect -224 -18806 -204 -12784
rect -140 -18806 -120 -12784
rect 3107 -12835 3211 -12437
rect 6386 -12488 6406 -6466
rect 6470 -12488 6490 -6466
rect 9717 -6517 9821 -6119
rect 12996 -6170 13016 -148
rect 13080 -6170 13100 -148
rect 16327 -199 16431 199
rect 19606 148 19626 6170
rect 19690 148 19710 6170
rect 19606 -148 19710 148
rect 13419 -200 19339 -199
rect 13419 -6118 13420 -200
rect 19338 -6118 19339 -200
rect 13419 -6119 19339 -6118
rect 12996 -6466 13100 -6170
rect 6809 -6518 12729 -6517
rect 6809 -12436 6810 -6518
rect 12728 -12436 12729 -6518
rect 6809 -12437 12729 -12436
rect 6386 -12784 6490 -12488
rect 199 -12836 6119 -12835
rect 199 -18754 200 -12836
rect 6118 -18754 6119 -12836
rect 199 -18755 6119 -18754
rect -224 -18954 -120 -18806
rect 3107 -18954 3211 -18755
rect 6386 -18806 6406 -12784
rect 6470 -18806 6490 -12784
rect 9717 -12835 9821 -12437
rect 12996 -12488 13016 -6466
rect 13080 -12488 13100 -6466
rect 16327 -6517 16431 -6119
rect 19606 -6170 19626 -148
rect 19690 -6170 19710 -148
rect 19606 -6466 19710 -6170
rect 13419 -6518 19339 -6517
rect 13419 -12436 13420 -6518
rect 19338 -12436 19339 -6518
rect 13419 -12437 19339 -12436
rect 12996 -12784 13100 -12488
rect 6809 -12836 12729 -12835
rect 6809 -18754 6810 -12836
rect 12728 -18754 12729 -12836
rect 6809 -18755 12729 -18754
rect 6386 -18954 6490 -18806
rect 9717 -18954 9821 -18755
rect 12996 -18806 13016 -12784
rect 13080 -18806 13100 -12784
rect 16327 -12835 16431 -12437
rect 19606 -12488 19626 -6466
rect 19690 -12488 19710 -6466
rect 19606 -12784 19710 -12488
rect 13419 -12836 19339 -12835
rect 13419 -18754 13420 -12836
rect 19338 -18754 19339 -12836
rect 13419 -18755 19339 -18754
rect 12996 -18954 13100 -18806
rect 16327 -18954 16431 -18755
rect 19606 -18806 19626 -12784
rect 19690 -18806 19710 -12784
rect 19606 -18954 19710 -18806
<< properties >>
string FIXED_BBOX 13340 12756 19418 18834
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 29.993 l 29.993 val 1.821k carea 2.00 cperi 0.19 nx 6 ny 6 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1702109072
<< metal3 >>
rect -16410 15652 -10038 15680
rect -16410 9628 -10122 15652
rect -10058 9628 -10038 15652
rect -16410 9600 -10038 9628
rect -9798 15652 -3426 15680
rect -9798 9628 -3510 15652
rect -3446 9628 -3426 15652
rect -9798 9600 -3426 9628
rect -3186 15652 3186 15680
rect -3186 9628 3102 15652
rect 3166 9628 3186 15652
rect -3186 9600 3186 9628
rect 3426 15652 9798 15680
rect 3426 9628 9714 15652
rect 9778 9628 9798 15652
rect 3426 9600 9798 9628
rect 10038 15652 16410 15680
rect 10038 9628 16326 15652
rect 16390 9628 16410 15652
rect 10038 9600 16410 9628
rect -16410 9332 -10038 9360
rect -16410 3308 -10122 9332
rect -10058 3308 -10038 9332
rect -16410 3280 -10038 3308
rect -9798 9332 -3426 9360
rect -9798 3308 -3510 9332
rect -3446 3308 -3426 9332
rect -9798 3280 -3426 3308
rect -3186 9332 3186 9360
rect -3186 3308 3102 9332
rect 3166 3308 3186 9332
rect -3186 3280 3186 3308
rect 3426 9332 9798 9360
rect 3426 3308 9714 9332
rect 9778 3308 9798 9332
rect 3426 3280 9798 3308
rect 10038 9332 16410 9360
rect 10038 3308 16326 9332
rect 16390 3308 16410 9332
rect 10038 3280 16410 3308
rect -16410 3012 -10038 3040
rect -16410 -3012 -10122 3012
rect -10058 -3012 -10038 3012
rect -16410 -3040 -10038 -3012
rect -9798 3012 -3426 3040
rect -9798 -3012 -3510 3012
rect -3446 -3012 -3426 3012
rect -9798 -3040 -3426 -3012
rect -3186 3012 3186 3040
rect -3186 -3012 3102 3012
rect 3166 -3012 3186 3012
rect -3186 -3040 3186 -3012
rect 3426 3012 9798 3040
rect 3426 -3012 9714 3012
rect 9778 -3012 9798 3012
rect 3426 -3040 9798 -3012
rect 10038 3012 16410 3040
rect 10038 -3012 16326 3012
rect 16390 -3012 16410 3012
rect 10038 -3040 16410 -3012
rect -16410 -3308 -10038 -3280
rect -16410 -9332 -10122 -3308
rect -10058 -9332 -10038 -3308
rect -16410 -9360 -10038 -9332
rect -9798 -3308 -3426 -3280
rect -9798 -9332 -3510 -3308
rect -3446 -9332 -3426 -3308
rect -9798 -9360 -3426 -9332
rect -3186 -3308 3186 -3280
rect -3186 -9332 3102 -3308
rect 3166 -9332 3186 -3308
rect -3186 -9360 3186 -9332
rect 3426 -3308 9798 -3280
rect 3426 -9332 9714 -3308
rect 9778 -9332 9798 -3308
rect 3426 -9360 9798 -9332
rect 10038 -3308 16410 -3280
rect 10038 -9332 16326 -3308
rect 16390 -9332 16410 -3308
rect 10038 -9360 16410 -9332
rect -16410 -9628 -10038 -9600
rect -16410 -15652 -10122 -9628
rect -10058 -15652 -10038 -9628
rect -16410 -15680 -10038 -15652
rect -9798 -9628 -3426 -9600
rect -9798 -15652 -3510 -9628
rect -3446 -15652 -3426 -9628
rect -9798 -15680 -3426 -15652
rect -3186 -9628 3186 -9600
rect -3186 -15652 3102 -9628
rect 3166 -15652 3186 -9628
rect -3186 -15680 3186 -15652
rect 3426 -9628 9798 -9600
rect 3426 -15652 9714 -9628
rect 9778 -15652 9798 -9628
rect 3426 -15680 9798 -15652
rect 10038 -9628 16410 -9600
rect 10038 -15652 16326 -9628
rect 16390 -15652 16410 -9628
rect 10038 -15680 16410 -15652
<< via3 >>
rect -10122 9628 -10058 15652
rect -3510 9628 -3446 15652
rect 3102 9628 3166 15652
rect 9714 9628 9778 15652
rect 16326 9628 16390 15652
rect -10122 3308 -10058 9332
rect -3510 3308 -3446 9332
rect 3102 3308 3166 9332
rect 9714 3308 9778 9332
rect 16326 3308 16390 9332
rect -10122 -3012 -10058 3012
rect -3510 -3012 -3446 3012
rect 3102 -3012 3166 3012
rect 9714 -3012 9778 3012
rect 16326 -3012 16390 3012
rect -10122 -9332 -10058 -3308
rect -3510 -9332 -3446 -3308
rect 3102 -9332 3166 -3308
rect 9714 -9332 9778 -3308
rect 16326 -9332 16390 -3308
rect -10122 -15652 -10058 -9628
rect -3510 -15652 -3446 -9628
rect 3102 -15652 3166 -9628
rect 9714 -15652 9778 -9628
rect 16326 -15652 16390 -9628
<< mimcap >>
rect -16370 15600 -10370 15640
rect -16370 9680 -16330 15600
rect -10410 9680 -10370 15600
rect -16370 9640 -10370 9680
rect -9758 15600 -3758 15640
rect -9758 9680 -9718 15600
rect -3798 9680 -3758 15600
rect -9758 9640 -3758 9680
rect -3146 15600 2854 15640
rect -3146 9680 -3106 15600
rect 2814 9680 2854 15600
rect -3146 9640 2854 9680
rect 3466 15600 9466 15640
rect 3466 9680 3506 15600
rect 9426 9680 9466 15600
rect 3466 9640 9466 9680
rect 10078 15600 16078 15640
rect 10078 9680 10118 15600
rect 16038 9680 16078 15600
rect 10078 9640 16078 9680
rect -16370 9280 -10370 9320
rect -16370 3360 -16330 9280
rect -10410 3360 -10370 9280
rect -16370 3320 -10370 3360
rect -9758 9280 -3758 9320
rect -9758 3360 -9718 9280
rect -3798 3360 -3758 9280
rect -9758 3320 -3758 3360
rect -3146 9280 2854 9320
rect -3146 3360 -3106 9280
rect 2814 3360 2854 9280
rect -3146 3320 2854 3360
rect 3466 9280 9466 9320
rect 3466 3360 3506 9280
rect 9426 3360 9466 9280
rect 3466 3320 9466 3360
rect 10078 9280 16078 9320
rect 10078 3360 10118 9280
rect 16038 3360 16078 9280
rect 10078 3320 16078 3360
rect -16370 2960 -10370 3000
rect -16370 -2960 -16330 2960
rect -10410 -2960 -10370 2960
rect -16370 -3000 -10370 -2960
rect -9758 2960 -3758 3000
rect -9758 -2960 -9718 2960
rect -3798 -2960 -3758 2960
rect -9758 -3000 -3758 -2960
rect -3146 2960 2854 3000
rect -3146 -2960 -3106 2960
rect 2814 -2960 2854 2960
rect -3146 -3000 2854 -2960
rect 3466 2960 9466 3000
rect 3466 -2960 3506 2960
rect 9426 -2960 9466 2960
rect 3466 -3000 9466 -2960
rect 10078 2960 16078 3000
rect 10078 -2960 10118 2960
rect 16038 -2960 16078 2960
rect 10078 -3000 16078 -2960
rect -16370 -3360 -10370 -3320
rect -16370 -9280 -16330 -3360
rect -10410 -9280 -10370 -3360
rect -16370 -9320 -10370 -9280
rect -9758 -3360 -3758 -3320
rect -9758 -9280 -9718 -3360
rect -3798 -9280 -3758 -3360
rect -9758 -9320 -3758 -9280
rect -3146 -3360 2854 -3320
rect -3146 -9280 -3106 -3360
rect 2814 -9280 2854 -3360
rect -3146 -9320 2854 -9280
rect 3466 -3360 9466 -3320
rect 3466 -9280 3506 -3360
rect 9426 -9280 9466 -3360
rect 3466 -9320 9466 -9280
rect 10078 -3360 16078 -3320
rect 10078 -9280 10118 -3360
rect 16038 -9280 16078 -3360
rect 10078 -9320 16078 -9280
rect -16370 -9680 -10370 -9640
rect -16370 -15600 -16330 -9680
rect -10410 -15600 -10370 -9680
rect -16370 -15640 -10370 -15600
rect -9758 -9680 -3758 -9640
rect -9758 -15600 -9718 -9680
rect -3798 -15600 -3758 -9680
rect -9758 -15640 -3758 -15600
rect -3146 -9680 2854 -9640
rect -3146 -15600 -3106 -9680
rect 2814 -15600 2854 -9680
rect -3146 -15640 2854 -15600
rect 3466 -9680 9466 -9640
rect 3466 -15600 3506 -9680
rect 9426 -15600 9466 -9680
rect 3466 -15640 9466 -15600
rect 10078 -9680 16078 -9640
rect 10078 -15600 10118 -9680
rect 16038 -15600 16078 -9680
rect 10078 -15640 16078 -15600
<< mimcapcontact >>
rect -16330 9680 -10410 15600
rect -9718 9680 -3798 15600
rect -3106 9680 2814 15600
rect 3506 9680 9426 15600
rect 10118 9680 16038 15600
rect -16330 3360 -10410 9280
rect -9718 3360 -3798 9280
rect -3106 3360 2814 9280
rect 3506 3360 9426 9280
rect 10118 3360 16038 9280
rect -16330 -2960 -10410 2960
rect -9718 -2960 -3798 2960
rect -3106 -2960 2814 2960
rect 3506 -2960 9426 2960
rect 10118 -2960 16038 2960
rect -16330 -9280 -10410 -3360
rect -9718 -9280 -3798 -3360
rect -3106 -9280 2814 -3360
rect 3506 -9280 9426 -3360
rect 10118 -9280 16038 -3360
rect -16330 -15600 -10410 -9680
rect -9718 -15600 -3798 -9680
rect -3106 -15600 2814 -9680
rect 3506 -15600 9426 -9680
rect 10118 -15600 16038 -9680
<< metal4 >>
rect -13422 15601 -13318 15800
rect -10142 15652 -10038 15800
rect -16331 15600 -10409 15601
rect -16331 9680 -16330 15600
rect -10410 9680 -10409 15600
rect -16331 9679 -10409 9680
rect -13422 9281 -13318 9679
rect -10142 9628 -10122 15652
rect -10058 9628 -10038 15652
rect -6810 15601 -6706 15800
rect -3530 15652 -3426 15800
rect -9719 15600 -3797 15601
rect -9719 9680 -9718 15600
rect -3798 9680 -3797 15600
rect -9719 9679 -3797 9680
rect -10142 9332 -10038 9628
rect -16331 9280 -10409 9281
rect -16331 3360 -16330 9280
rect -10410 3360 -10409 9280
rect -16331 3359 -10409 3360
rect -13422 2961 -13318 3359
rect -10142 3308 -10122 9332
rect -10058 3308 -10038 9332
rect -6810 9281 -6706 9679
rect -3530 9628 -3510 15652
rect -3446 9628 -3426 15652
rect -198 15601 -94 15800
rect 3082 15652 3186 15800
rect -3107 15600 2815 15601
rect -3107 9680 -3106 15600
rect 2814 9680 2815 15600
rect -3107 9679 2815 9680
rect -3530 9332 -3426 9628
rect -9719 9280 -3797 9281
rect -9719 3360 -9718 9280
rect -3798 3360 -3797 9280
rect -9719 3359 -3797 3360
rect -10142 3012 -10038 3308
rect -16331 2960 -10409 2961
rect -16331 -2960 -16330 2960
rect -10410 -2960 -10409 2960
rect -16331 -2961 -10409 -2960
rect -13422 -3359 -13318 -2961
rect -10142 -3012 -10122 3012
rect -10058 -3012 -10038 3012
rect -6810 2961 -6706 3359
rect -3530 3308 -3510 9332
rect -3446 3308 -3426 9332
rect -198 9281 -94 9679
rect 3082 9628 3102 15652
rect 3166 9628 3186 15652
rect 6414 15601 6518 15800
rect 9694 15652 9798 15800
rect 3505 15600 9427 15601
rect 3505 9680 3506 15600
rect 9426 9680 9427 15600
rect 3505 9679 9427 9680
rect 3082 9332 3186 9628
rect -3107 9280 2815 9281
rect -3107 3360 -3106 9280
rect 2814 3360 2815 9280
rect -3107 3359 2815 3360
rect -3530 3012 -3426 3308
rect -9719 2960 -3797 2961
rect -9719 -2960 -9718 2960
rect -3798 -2960 -3797 2960
rect -9719 -2961 -3797 -2960
rect -10142 -3308 -10038 -3012
rect -16331 -3360 -10409 -3359
rect -16331 -9280 -16330 -3360
rect -10410 -9280 -10409 -3360
rect -16331 -9281 -10409 -9280
rect -13422 -9679 -13318 -9281
rect -10142 -9332 -10122 -3308
rect -10058 -9332 -10038 -3308
rect -6810 -3359 -6706 -2961
rect -3530 -3012 -3510 3012
rect -3446 -3012 -3426 3012
rect -198 2961 -94 3359
rect 3082 3308 3102 9332
rect 3166 3308 3186 9332
rect 6414 9281 6518 9679
rect 9694 9628 9714 15652
rect 9778 9628 9798 15652
rect 13026 15601 13130 15800
rect 16306 15652 16410 15800
rect 10117 15600 16039 15601
rect 10117 9680 10118 15600
rect 16038 9680 16039 15600
rect 10117 9679 16039 9680
rect 9694 9332 9798 9628
rect 3505 9280 9427 9281
rect 3505 3360 3506 9280
rect 9426 3360 9427 9280
rect 3505 3359 9427 3360
rect 3082 3012 3186 3308
rect -3107 2960 2815 2961
rect -3107 -2960 -3106 2960
rect 2814 -2960 2815 2960
rect -3107 -2961 2815 -2960
rect -3530 -3308 -3426 -3012
rect -9719 -3360 -3797 -3359
rect -9719 -9280 -9718 -3360
rect -3798 -9280 -3797 -3360
rect -9719 -9281 -3797 -9280
rect -10142 -9628 -10038 -9332
rect -16331 -9680 -10409 -9679
rect -16331 -15600 -16330 -9680
rect -10410 -15600 -10409 -9680
rect -16331 -15601 -10409 -15600
rect -13422 -15800 -13318 -15601
rect -10142 -15652 -10122 -9628
rect -10058 -15652 -10038 -9628
rect -6810 -9679 -6706 -9281
rect -3530 -9332 -3510 -3308
rect -3446 -9332 -3426 -3308
rect -198 -3359 -94 -2961
rect 3082 -3012 3102 3012
rect 3166 -3012 3186 3012
rect 6414 2961 6518 3359
rect 9694 3308 9714 9332
rect 9778 3308 9798 9332
rect 13026 9281 13130 9679
rect 16306 9628 16326 15652
rect 16390 9628 16410 15652
rect 16306 9332 16410 9628
rect 10117 9280 16039 9281
rect 10117 3360 10118 9280
rect 16038 3360 16039 9280
rect 10117 3359 16039 3360
rect 9694 3012 9798 3308
rect 3505 2960 9427 2961
rect 3505 -2960 3506 2960
rect 9426 -2960 9427 2960
rect 3505 -2961 9427 -2960
rect 3082 -3308 3186 -3012
rect -3107 -3360 2815 -3359
rect -3107 -9280 -3106 -3360
rect 2814 -9280 2815 -3360
rect -3107 -9281 2815 -9280
rect -3530 -9628 -3426 -9332
rect -9719 -9680 -3797 -9679
rect -9719 -15600 -9718 -9680
rect -3798 -15600 -3797 -9680
rect -9719 -15601 -3797 -15600
rect -10142 -15800 -10038 -15652
rect -6810 -15800 -6706 -15601
rect -3530 -15652 -3510 -9628
rect -3446 -15652 -3426 -9628
rect -198 -9679 -94 -9281
rect 3082 -9332 3102 -3308
rect 3166 -9332 3186 -3308
rect 6414 -3359 6518 -2961
rect 9694 -3012 9714 3012
rect 9778 -3012 9798 3012
rect 13026 2961 13130 3359
rect 16306 3308 16326 9332
rect 16390 3308 16410 9332
rect 16306 3012 16410 3308
rect 10117 2960 16039 2961
rect 10117 -2960 10118 2960
rect 16038 -2960 16039 2960
rect 10117 -2961 16039 -2960
rect 9694 -3308 9798 -3012
rect 3505 -3360 9427 -3359
rect 3505 -9280 3506 -3360
rect 9426 -9280 9427 -3360
rect 3505 -9281 9427 -9280
rect 3082 -9628 3186 -9332
rect -3107 -9680 2815 -9679
rect -3107 -15600 -3106 -9680
rect 2814 -15600 2815 -9680
rect -3107 -15601 2815 -15600
rect -3530 -15800 -3426 -15652
rect -198 -15800 -94 -15601
rect 3082 -15652 3102 -9628
rect 3166 -15652 3186 -9628
rect 6414 -9679 6518 -9281
rect 9694 -9332 9714 -3308
rect 9778 -9332 9798 -3308
rect 13026 -3359 13130 -2961
rect 16306 -3012 16326 3012
rect 16390 -3012 16410 3012
rect 16306 -3308 16410 -3012
rect 10117 -3360 16039 -3359
rect 10117 -9280 10118 -3360
rect 16038 -9280 16039 -3360
rect 10117 -9281 16039 -9280
rect 9694 -9628 9798 -9332
rect 3505 -9680 9427 -9679
rect 3505 -15600 3506 -9680
rect 9426 -15600 9427 -9680
rect 3505 -15601 9427 -15600
rect 3082 -15800 3186 -15652
rect 6414 -15800 6518 -15601
rect 9694 -15652 9714 -9628
rect 9778 -15652 9798 -9628
rect 13026 -9679 13130 -9281
rect 16306 -9332 16326 -3308
rect 16390 -9332 16410 -3308
rect 16306 -9628 16410 -9332
rect 10117 -9680 16039 -9679
rect 10117 -15600 10118 -9680
rect 16038 -15600 16039 -9680
rect 10117 -15601 16039 -15600
rect 9694 -15800 9798 -15652
rect 13026 -15800 13130 -15601
rect 16306 -15652 16326 -9628
rect 16390 -15652 16410 -9628
rect 16306 -15800 16410 -15652
<< properties >>
string FIXED_BBOX 10038 9600 16118 15680
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 5 ny 5 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

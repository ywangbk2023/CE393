magic
tech sky130A
magscale 1 2
timestamp 1702109646
<< nwell >>
rect 1458 2484 2236 2508
rect 338 1626 2344 2484
rect -408 1474 3350 1626
rect -410 1118 3356 1474
rect -410 1108 576 1118
rect 594 1108 638 1110
rect 658 1108 3356 1118
rect -410 1106 3356 1108
rect 594 1048 638 1106
rect 1972 1040 2006 1106
rect 42 264 88 272
rect 1748 268 1794 274
rect -40 134 -38 168
rect 10 104 342 264
rect 1746 204 1798 268
rect 1800 236 1960 254
rect 18 -524 330 104
rect 692 -76 3044 204
rect 1706 -80 2036 -76
rect 16 -602 346 -524
rect 470 -602 538 -524
rect 1724 -802 2036 -80
rect 732 -2488 1610 -2448
rect 1790 -2488 2668 -2448
rect 2798 -2488 3676 -2448
rect 1650 -2516 1752 -2506
rect 614 -2522 648 -2516
rect 1622 -2522 1778 -2516
rect 2752 -2522 2786 -2516
rect 1650 -2698 1754 -2522
rect 1650 -2710 1752 -2698
rect 2360 -4294 2610 -4276
rect 1724 -4316 2610 -4294
rect 604 -5172 2610 -4316
<< pmos >>
rect 470 -540 538 -524
<< ndiff >>
rect 2274 -1604 2284 -1570
rect 1474 -1680 1486 -1666
rect 2842 -1684 2844 -1496
<< pdiff >>
rect 1650 -2698 1754 -2522
<< poly >>
rect 1458 2498 2236 2508
rect 1458 2496 2128 2498
rect 1458 2462 1646 2496
rect 1680 2462 1796 2496
rect 1830 2462 1966 2496
rect 2000 2464 2128 2496
rect 2164 2464 2236 2498
rect 2000 2462 2236 2464
rect 1458 2450 2236 2462
rect 1458 2432 2190 2450
rect 458 2118 558 2206
rect 616 2118 716 2206
rect 774 2118 874 2206
rect 932 2118 1032 2206
rect 1090 2118 1190 2206
rect 458 2058 480 2118
rect 534 2058 636 2118
rect 690 2116 956 2118
rect 690 2058 798 2116
rect 458 1966 558 2058
rect 616 1966 716 2058
rect 774 2056 798 2058
rect 852 2058 956 2116
rect 1010 2116 1190 2118
rect 1010 2058 1108 2116
rect 852 2056 874 2058
rect 774 1966 874 2056
rect 932 1966 1032 2058
rect 1090 2056 1108 2058
rect 1162 2056 1190 2116
rect 1090 1966 1190 2056
rect 1456 1716 2190 1746
rect 1456 1714 1806 1716
rect 1456 1672 1488 1714
rect 1526 1672 1648 1714
rect 1686 1674 1806 1714
rect 1844 1714 2118 1716
rect 1844 1674 1962 1714
rect 1686 1672 1962 1674
rect 2000 1674 2118 1714
rect 2156 1674 2190 1716
rect 2000 1672 2190 1674
rect 1456 1662 2190 1672
rect 94 -142 254 246
rect 94 -216 140 -142
rect 204 -216 254 -142
rect 94 -232 254 -216
rect 1800 -140 1960 254
rect 1800 -214 1846 -140
rect 1910 -214 1960 -140
rect 1800 -230 1960 -214
rect -184 -622 -136 -524
rect 470 -566 538 -540
rect 480 -622 528 -566
rect -194 -630 -126 -622
rect -194 -698 -178 -630
rect -142 -698 -126 -630
rect -194 -708 -126 -698
rect 470 -630 538 -622
rect 470 -698 486 -630
rect 522 -698 538 -630
rect 470 -708 538 -698
rect -76 -750 -8 -740
rect -124 -818 -60 -750
rect -24 -818 -8 -750
rect -124 -828 -8 -818
rect 356 -750 424 -740
rect 356 -818 372 -750
rect 408 -818 472 -750
rect 972 -756 1172 -708
rect 1230 -756 1430 -704
rect 356 -828 472 -818
rect 770 -762 1430 -756
rect 2330 -758 2530 -702
rect 2588 -758 2788 -696
rect 770 -818 1788 -762
rect 2330 -766 2788 -758
rect 770 -824 1694 -818
rect -124 -870 -76 -828
rect 424 -870 472 -828
rect 972 -830 1430 -824
rect 972 -870 1172 -830
rect 1230 -870 1430 -830
rect 1678 -894 1694 -824
rect 1772 -894 1788 -818
rect 1678 -910 1788 -894
rect 1964 -818 2990 -766
rect 1964 -894 1980 -818
rect 2058 -828 2990 -818
rect 2058 -894 2074 -828
rect 2330 -832 2788 -828
rect 2330 -862 2530 -832
rect 2588 -856 2788 -832
rect 1964 -910 2074 -894
rect 1820 -1240 1980 -1216
rect 1820 -1352 1848 -1240
rect 1948 -1352 1980 -1240
rect 1820 -1386 1980 -1352
rect 1818 -1640 1980 -1386
rect 1820 -1670 1980 -1640
rect -276 -2420 602 -2410
rect -276 -2446 -192 -2420
rect -230 -2460 -192 -2446
rect -150 -2422 166 -2420
rect -150 -2460 -18 -2422
rect -230 -2462 -18 -2460
rect 24 -2460 166 -2422
rect 208 -2460 322 -2420
rect 364 -2460 602 -2420
rect 732 -2420 1610 -2410
rect 732 -2446 816 -2420
rect 24 -2462 602 -2460
rect -230 -2488 602 -2462
rect 778 -2460 816 -2446
rect 858 -2422 1174 -2420
rect 858 -2460 990 -2422
rect 778 -2462 990 -2460
rect 1032 -2460 1174 -2422
rect 1216 -2460 1330 -2420
rect 1372 -2460 1610 -2420
rect 1032 -2462 1610 -2460
rect 778 -2488 1610 -2462
rect 1790 -2420 2668 -2410
rect 1790 -2460 2028 -2420
rect 2070 -2460 2184 -2420
rect 2226 -2422 2542 -2420
rect 2226 -2460 2368 -2422
rect 1790 -2462 2368 -2460
rect 2410 -2460 2542 -2422
rect 2584 -2446 2668 -2420
rect 2798 -2420 3676 -2410
rect 2584 -2460 2622 -2446
rect 2410 -2462 2622 -2460
rect 1790 -2488 2622 -2462
rect 2798 -2460 3036 -2420
rect 3078 -2460 3192 -2420
rect 3234 -2422 3550 -2420
rect 3234 -2460 3376 -2422
rect 2798 -2462 3376 -2460
rect 3418 -2460 3550 -2422
rect 3592 -2446 3676 -2420
rect 3592 -2460 3630 -2446
rect 3418 -2462 3630 -2460
rect 2798 -2488 3630 -2462
rect 2360 -4294 2440 -4276
rect 1724 -4302 2502 -4294
rect 1724 -4304 2394 -4302
rect 1724 -4338 1912 -4304
rect 1946 -4338 2062 -4304
rect 2096 -4338 2232 -4304
rect 2266 -4336 2394 -4304
rect 2430 -4336 2502 -4302
rect 2266 -4338 2502 -4336
rect 1724 -4350 2502 -4338
rect 1724 -4368 2456 -4350
rect 724 -4682 824 -4594
rect 882 -4682 982 -4594
rect 1040 -4682 1140 -4594
rect 1198 -4682 1298 -4594
rect 1356 -4682 1456 -4594
rect 724 -4742 746 -4682
rect 800 -4742 902 -4682
rect 956 -4684 1222 -4682
rect 956 -4742 1064 -4684
rect 724 -4834 824 -4742
rect 882 -4834 982 -4742
rect 1040 -4744 1064 -4742
rect 1118 -4742 1222 -4684
rect 1276 -4684 1456 -4682
rect 1276 -4742 1374 -4684
rect 1118 -4744 1140 -4742
rect 1040 -4834 1140 -4744
rect 1198 -4834 1298 -4742
rect 1356 -4744 1374 -4742
rect 1428 -4744 1456 -4684
rect 1356 -4834 1456 -4744
rect 1722 -5084 2456 -5054
rect 1722 -5086 2072 -5084
rect 1722 -5128 1754 -5086
rect 1792 -5128 1914 -5086
rect 1952 -5126 2072 -5086
rect 2110 -5086 2456 -5084
rect 2110 -5126 2228 -5086
rect 1952 -5128 2228 -5126
rect 2266 -5128 2456 -5086
rect 1722 -5138 2456 -5128
<< polycont >>
rect 1646 2462 1680 2496
rect 1796 2462 1830 2496
rect 1966 2462 2000 2496
rect 2128 2464 2164 2498
rect 480 2058 534 2118
rect 636 2058 690 2118
rect 798 2056 852 2116
rect 956 2058 1010 2118
rect 1108 2056 1162 2116
rect 1488 1672 1526 1714
rect 1648 1672 1686 1714
rect 1806 1674 1844 1716
rect 1962 1672 2000 1714
rect 2118 1674 2156 1716
rect 140 -216 204 -142
rect 1846 -214 1910 -140
rect -178 -698 -142 -630
rect 486 -698 522 -630
rect -60 -818 -24 -750
rect 372 -818 408 -750
rect 1694 -894 1772 -818
rect 1980 -894 2058 -818
rect 1848 -1352 1948 -1240
rect -192 -2460 -150 -2420
rect -18 -2462 24 -2422
rect 166 -2460 208 -2420
rect 322 -2460 364 -2420
rect 816 -2460 858 -2420
rect 990 -2462 1032 -2422
rect 1174 -2460 1216 -2420
rect 1330 -2460 1372 -2420
rect 2028 -2460 2070 -2420
rect 2184 -2460 2226 -2420
rect 2368 -2462 2410 -2422
rect 2542 -2460 2584 -2420
rect 3036 -2460 3078 -2420
rect 3192 -2460 3234 -2420
rect 3376 -2462 3418 -2422
rect 3550 -2460 3592 -2420
rect 1912 -4338 1946 -4304
rect 2062 -4338 2096 -4304
rect 2232 -4338 2266 -4304
rect 2394 -4336 2430 -4302
rect 746 -4742 800 -4682
rect 902 -4742 956 -4682
rect 1064 -4744 1118 -4684
rect 1222 -4742 1276 -4682
rect 1374 -4744 1428 -4684
rect 1754 -5128 1792 -5086
rect 1914 -5128 1952 -5086
rect 2072 -5126 2110 -5084
rect 2228 -5128 2266 -5086
<< locali >>
rect 2162 2702 2248 2770
rect 2170 2508 2238 2702
rect 1570 2498 2238 2508
rect 1570 2496 2128 2498
rect 412 2450 1446 2484
rect 412 2390 446 2450
rect 728 2400 762 2450
rect 1044 2448 1446 2450
rect 1044 2402 1078 2448
rect 1412 2408 1446 2448
rect 1570 2462 1646 2496
rect 1680 2462 1796 2496
rect 1830 2462 1966 2496
rect 2000 2464 2128 2496
rect 2164 2464 2238 2498
rect 2000 2462 2238 2464
rect 1570 2450 2238 2462
rect 1570 2402 1604 2450
rect 1886 2400 1920 2450
rect 2170 2448 2238 2450
rect 2202 2390 2236 2448
rect 570 2154 606 2216
rect 886 2154 920 2214
rect 1202 2154 1236 2206
rect 412 2118 1236 2154
rect 1412 2154 1446 2206
rect 1728 2154 1762 2214
rect 2042 2154 2078 2216
rect 1412 2120 2078 2154
rect 412 2058 480 2118
rect 534 2058 636 2118
rect 690 2116 956 2118
rect 690 2058 798 2116
rect 412 2056 798 2058
rect 852 2058 956 2116
rect 1010 2116 1236 2118
rect 1010 2058 1108 2116
rect 852 2056 1108 2058
rect 1162 2056 1236 2116
rect 412 2008 1236 2056
rect 1568 2010 2236 2044
rect 412 1950 446 2008
rect 728 1960 762 2008
rect 1044 1962 1078 2008
rect 1570 1962 1604 2010
rect 1886 1960 1920 2010
rect 2202 1950 2236 2010
rect 570 1714 606 1776
rect 886 1714 920 1774
rect 1202 1714 1236 1766
rect 1412 1728 1446 1766
rect 1728 1728 1762 1774
rect 2042 1728 2078 1776
rect 1412 1718 2190 1728
rect 1412 1716 2110 1718
rect 1412 1714 1806 1716
rect 570 1680 1488 1714
rect 1456 1672 1488 1680
rect 1526 1672 1648 1714
rect 1686 1674 1806 1714
rect 1844 1714 2110 1716
rect 1844 1674 1962 1714
rect 1686 1672 1962 1674
rect 2000 1672 2110 1714
rect 2158 1672 2190 1718
rect 1456 1662 2190 1672
rect -346 1306 -126 1368
rect -346 1188 -302 1306
rect -174 1188 -126 1306
rect -346 1118 -126 1188
rect 258 1352 308 1368
rect 258 1126 266 1352
rect 300 1126 308 1352
rect 258 1118 308 1126
rect 1960 1360 2022 1368
rect 1960 1124 1972 1360
rect 2006 1124 2022 1360
rect 1960 1118 2022 1124
rect 266 1042 300 1118
rect 1972 1040 2006 1118
rect -40 134 -38 168
rect 94 -138 254 -120
rect 94 -220 136 -138
rect 208 -220 254 -138
rect 94 -232 254 -220
rect 1800 -136 1960 -118
rect 1800 -218 1842 -136
rect 1914 -218 1960 -136
rect 1800 -230 1960 -218
rect -282 -756 -248 -544
rect -194 -630 -126 -622
rect -194 -698 -178 -630
rect -142 -698 -126 -630
rect -194 -708 -126 -698
rect 470 -630 538 -622
rect 470 -698 486 -630
rect 522 -698 538 -630
rect 470 -708 538 -698
rect -76 -750 -8 -740
rect 356 -750 424 -740
rect 596 -750 630 -544
rect -298 -762 -232 -756
rect -298 -826 -282 -762
rect -248 -826 -232 -762
rect -298 -832 -232 -826
rect -76 -818 -60 -750
rect -24 -818 372 -750
rect 408 -818 630 -750
rect 1184 -784 1218 -744
rect -76 -828 -8 -818
rect 356 -828 424 -818
rect -282 -872 -248 -832
rect 596 -872 630 -818
rect 770 -826 1606 -784
rect 2542 -790 2576 -744
rect 770 -1226 812 -826
rect 1184 -876 1218 -826
rect 1184 -902 1218 -884
rect 1564 -982 1606 -826
rect 1678 -818 1788 -790
rect 1678 -894 1694 -818
rect 1772 -894 1788 -818
rect 1678 -910 1788 -894
rect 1964 -818 2074 -802
rect 1964 -894 1980 -818
rect 2058 -894 2074 -818
rect 2542 -832 3016 -790
rect 2542 -876 2576 -832
rect 1964 -910 2074 -894
rect 2974 -936 3016 -832
rect 2964 -942 3026 -936
rect 1554 -988 1616 -982
rect 1554 -1032 1568 -988
rect 1604 -1032 1616 -988
rect 2964 -986 2978 -942
rect 3014 -986 3026 -942
rect 2964 -992 3026 -986
rect 1554 -1038 1616 -1032
rect 756 -1238 826 -1226
rect 756 -1280 772 -1238
rect 810 -1280 826 -1238
rect 756 -1294 826 -1280
rect 1820 -1234 1980 -1216
rect 1820 -1362 1842 -1234
rect 1956 -1362 1980 -1234
rect 1820 -1374 1980 -1362
rect 1774 -1600 2300 -1552
rect 1774 -1668 1808 -1600
rect 2284 -1604 2286 -1600
rect -64 -2118 -30 -2072
rect 378 -2118 412 -2072
rect 1466 -2074 1782 -2026
rect 1992 -2118 2026 -1658
rect -326 -2124 -22 -2118
rect -326 -2162 -64 -2124
rect -326 -2322 -266 -2162
rect -126 -2322 -64 -2162
rect -326 -2360 -64 -2322
rect -30 -2360 -22 -2124
rect -326 -2368 -22 -2360
rect 370 -2124 420 -2118
rect 370 -2360 378 -2124
rect 412 -2360 420 -2124
rect 370 -2368 420 -2360
rect 1984 -2124 2034 -2118
rect 1984 -2360 1992 -2124
rect 2026 -2360 2034 -2124
rect 1984 -2368 2034 -2360
rect -276 -2418 602 -2410
rect -276 -2420 530 -2418
rect -276 -2460 -192 -2420
rect -150 -2422 166 -2420
rect -150 -2460 -18 -2422
rect -276 -2462 -18 -2460
rect 24 -2460 166 -2422
rect 208 -2460 322 -2420
rect 364 -2460 530 -2420
rect 24 -2462 530 -2460
rect 566 -2462 602 -2418
rect -276 -2470 602 -2462
rect 732 -2420 1478 -2410
rect 732 -2460 816 -2420
rect 858 -2422 1174 -2420
rect 858 -2460 990 -2422
rect 732 -2462 990 -2460
rect 1032 -2460 1174 -2422
rect 1216 -2460 1330 -2420
rect 1372 -2460 1478 -2420
rect 1032 -2462 1478 -2460
rect 732 -2470 1478 -2462
rect -276 -2506 -242 -2470
rect 80 -2532 114 -2470
rect 436 -2530 470 -2470
rect 732 -2506 766 -2470
rect 1088 -2532 1122 -2470
rect 1444 -2530 1478 -2470
rect 1922 -2420 2668 -2410
rect 1922 -2460 2028 -2420
rect 2070 -2460 2184 -2420
rect 2226 -2422 2542 -2420
rect 2226 -2460 2368 -2422
rect 1922 -2462 2368 -2460
rect 2410 -2460 2542 -2422
rect 2584 -2460 2668 -2420
rect 2410 -2462 2668 -2460
rect 1922 -2470 2668 -2462
rect 2798 -2418 3676 -2410
rect 2798 -2462 2832 -2418
rect 2890 -2420 3676 -2418
rect 2890 -2460 3036 -2420
rect 3078 -2460 3192 -2420
rect 3234 -2422 3550 -2420
rect 3234 -2460 3376 -2422
rect 2890 -2462 3376 -2460
rect 3418 -2460 3550 -2422
rect 3592 -2460 3676 -2420
rect 3418 -2462 3676 -2460
rect 2798 -2470 3676 -2462
rect 1650 -2522 1752 -2506
rect -98 -2780 -64 -2596
rect 258 -2780 292 -2710
rect 614 -2780 648 -2714
rect 732 -2780 766 -2712
rect -98 -2814 766 -2780
rect 910 -2780 944 -2596
rect 1650 -2698 1754 -2522
rect 1922 -2530 1956 -2470
rect 2278 -2532 2312 -2470
rect 2634 -2506 2668 -2470
rect 2930 -2530 2964 -2470
rect 3286 -2532 3320 -2470
rect 3642 -2506 3676 -2470
rect 1650 -2710 1752 -2698
rect 1266 -2780 1300 -2710
rect 1622 -2780 1656 -2714
rect 910 -2814 1656 -2780
rect 1744 -2780 1778 -2714
rect 2100 -2780 2134 -2710
rect 2456 -2780 2490 -2596
rect 1744 -2814 2490 -2780
rect 2634 -2780 2668 -2712
rect 2752 -2780 2786 -2714
rect 3108 -2780 3142 -2710
rect 3464 -2780 3498 -2596
rect 2634 -2814 3498 -2780
rect 2360 -4294 2440 -4276
rect 1836 -4304 2374 -4294
rect 2424 -4302 2502 -4294
rect 678 -4350 1712 -4316
rect 678 -4410 712 -4350
rect 994 -4400 1028 -4350
rect 1310 -4352 1712 -4350
rect 1310 -4398 1344 -4352
rect 1678 -4392 1712 -4352
rect 1836 -4338 1912 -4304
rect 1946 -4338 2062 -4304
rect 2096 -4338 2232 -4304
rect 2266 -4338 2374 -4304
rect 2430 -4336 2502 -4302
rect 1836 -4340 2374 -4338
rect 2424 -4340 2502 -4336
rect 1836 -4350 2502 -4340
rect 1836 -4398 1870 -4350
rect 2152 -4400 2186 -4350
rect 2468 -4410 2502 -4350
rect 836 -4646 872 -4584
rect 1152 -4646 1186 -4586
rect 1468 -4646 1502 -4594
rect 678 -4682 1502 -4646
rect 1678 -4646 1712 -4594
rect 1994 -4646 2028 -4586
rect 2308 -4646 2344 -4584
rect 1678 -4680 2344 -4646
rect 678 -4742 746 -4682
rect 800 -4742 902 -4682
rect 956 -4684 1222 -4682
rect 956 -4742 1064 -4684
rect 678 -4744 1064 -4742
rect 1118 -4742 1222 -4684
rect 1276 -4684 1502 -4682
rect 1276 -4742 1374 -4684
rect 1118 -4744 1374 -4742
rect 1428 -4744 1502 -4684
rect 678 -4792 1502 -4744
rect 1834 -4790 2502 -4756
rect 678 -4850 712 -4792
rect 994 -4840 1028 -4792
rect 1310 -4838 1344 -4792
rect 1836 -4838 1870 -4790
rect 2152 -4840 2186 -4790
rect 2468 -4850 2502 -4790
rect 836 -5086 872 -5024
rect 1152 -5086 1186 -5026
rect 1468 -5086 1502 -5034
rect 1678 -5072 1712 -5034
rect 1994 -5072 2028 -5026
rect 2308 -5070 2344 -5024
rect 2308 -5072 2456 -5070
rect 1678 -5084 2456 -5072
rect 1678 -5086 2072 -5084
rect 836 -5120 1754 -5086
rect 1722 -5128 1754 -5120
rect 1792 -5128 1914 -5086
rect 1952 -5126 2072 -5086
rect 2110 -5086 2456 -5084
rect 2110 -5126 2228 -5086
rect 1952 -5128 2228 -5126
rect 2266 -5128 2456 -5086
rect 1722 -5138 2456 -5128
<< viali >>
rect 2110 1716 2158 1718
rect 2110 1674 2118 1716
rect 2118 1674 2156 1716
rect 2156 1674 2158 1716
rect 2110 1672 2158 1674
rect -302 1188 -174 1306
rect 266 1126 300 1352
rect 1972 1124 2006 1360
rect 136 -142 208 -138
rect 136 -216 140 -142
rect 140 -216 204 -142
rect 204 -216 208 -142
rect 136 -220 208 -216
rect 1842 -140 1914 -136
rect 1842 -214 1846 -140
rect 1846 -214 1910 -140
rect 1910 -214 1914 -140
rect 1842 -218 1914 -214
rect -178 -682 -142 -648
rect -282 -826 -248 -762
rect 1568 -1032 1604 -988
rect 2978 -986 3014 -942
rect 772 -1280 810 -1238
rect 1842 -1240 1956 -1234
rect 1842 -1352 1848 -1240
rect 1848 -1352 1948 -1240
rect 1948 -1352 1956 -1240
rect 1842 -1362 1956 -1352
rect -266 -2322 -126 -2162
rect -64 -2360 -30 -2124
rect 378 -2360 412 -2124
rect 1992 -2360 2026 -2124
rect 530 -2462 566 -2418
rect 2832 -2462 2890 -2418
rect 2374 -4302 2424 -4294
rect 2374 -4336 2394 -4302
rect 2394 -4336 2424 -4302
rect 2374 -4340 2424 -4336
<< metal1 >>
rect 2162 2702 2248 2770
rect 2092 1722 2190 1728
rect 2092 1666 2108 1722
rect 2172 1666 2190 1722
rect 2092 1648 2190 1666
rect -346 1360 3250 1368
rect -346 1352 1972 1360
rect -346 1306 266 1352
rect -346 1188 -302 1306
rect -174 1188 266 1306
rect -346 1126 266 1188
rect 300 1126 1972 1352
rect -346 1124 1972 1126
rect 2006 1124 3250 1360
rect -346 1118 3250 1124
rect 42 216 88 272
rect -30 118 384 216
rect 1748 204 1794 274
rect 714 190 808 204
rect 714 -62 728 190
rect 784 -62 808 190
rect 714 -76 808 -62
rect 1590 198 1682 204
rect 1590 -66 1612 198
rect 1664 -66 1682 198
rect 1590 -76 1682 -66
rect 1732 198 1808 204
rect 1732 -70 1744 198
rect 1800 -70 1808 198
rect 1732 -76 1808 -70
rect 2056 196 2084 204
rect 2974 198 3064 212
rect 2056 -66 2064 196
rect 2056 -76 2084 -66
rect 2974 -72 2990 198
rect 3044 -72 3064 198
rect 2974 -88 3064 -72
rect 94 -134 254 -120
rect 94 -224 132 -134
rect 212 -224 254 -134
rect 94 -232 254 -224
rect 1800 -132 1960 -118
rect 1800 -222 1838 -132
rect 1918 -222 1960 -132
rect 1800 -230 1960 -222
rect -296 -648 -116 -642
rect -296 -682 -178 -648
rect -142 -682 -116 -648
rect -296 -690 -116 -682
rect -298 -762 -232 -756
rect -298 -826 -292 -762
rect -238 -826 -232 -762
rect -298 -832 -232 -826
rect 1678 -802 1788 -774
rect 1678 -904 1684 -802
rect 1782 -904 1788 -802
rect 1678 -910 1788 -904
rect 2954 -940 3038 -936
rect 1544 -982 1628 -980
rect 1544 -1034 1560 -982
rect 1614 -1034 1628 -982
rect 2954 -1002 2968 -940
rect 3022 -992 3038 -940
rect 3022 -1002 3034 -992
rect 2954 -1010 3034 -1002
rect 1544 -1040 1628 -1034
rect 756 -1236 826 -1226
rect 756 -1290 764 -1236
rect 820 -1290 826 -1236
rect 756 -1294 826 -1290
rect 1814 -1232 1986 -1216
rect 1814 -1366 1838 -1232
rect 1960 -1366 1986 -1232
rect 1814 -1374 1986 -1366
rect 2260 -1486 2322 -1450
rect 906 -1506 984 -1490
rect 906 -1682 914 -1506
rect 966 -1682 984 -1506
rect 906 -1694 984 -1682
rect 1418 -1512 1500 -1490
rect 1418 -1680 1432 -1512
rect 1486 -1680 1500 -1512
rect 2260 -1494 2336 -1486
rect 2260 -1612 2274 -1494
rect 1418 -1694 1500 -1680
rect 2268 -1682 2274 -1612
rect 2328 -1682 2336 -1494
rect 2268 -1690 2336 -1682
rect 2788 -1496 2860 -1486
rect 2788 -1684 2792 -1496
rect 2844 -1684 2860 -1496
rect 2788 -1690 2860 -1684
rect 1460 -1696 1500 -1694
rect -326 -2118 -82 -2116
rect -326 -2124 3294 -2118
rect -326 -2162 -64 -2124
rect -326 -2322 -266 -2162
rect -126 -2322 -64 -2162
rect -326 -2360 -64 -2322
rect -30 -2360 378 -2124
rect 412 -2360 1992 -2124
rect 2026 -2360 3294 -2124
rect -326 -2368 3294 -2360
rect 456 -2414 602 -2410
rect 456 -2466 522 -2414
rect 574 -2466 602 -2414
rect 456 -2470 602 -2466
rect 2798 -2414 2932 -2410
rect 2798 -2466 2828 -2414
rect 2894 -2466 2932 -2414
rect 2798 -2470 2932 -2466
rect 1616 -2710 1784 -2510
rect 1668 -2872 1732 -2710
rect 1658 -2882 1742 -2872
rect 1658 -2934 1674 -2882
rect 1726 -2934 1742 -2882
rect 1658 -2942 1742 -2934
rect 2360 -4290 2440 -4276
rect 2360 -4344 2368 -4290
rect 2430 -4344 2440 -4290
rect 2360 -4350 2440 -4344
rect 2368 -5140 2458 -5070
<< via1 >>
rect 2108 1718 2172 1722
rect 2108 1672 2110 1718
rect 2110 1672 2158 1718
rect 2158 1672 2172 1718
rect 2108 1666 2172 1672
rect 728 -62 784 190
rect 1612 -66 1664 198
rect 1744 -70 1800 198
rect 2064 -66 2124 196
rect 2990 -72 3044 198
rect 132 -138 212 -134
rect 132 -220 136 -138
rect 136 -220 208 -138
rect 208 -220 212 -138
rect 132 -224 212 -220
rect 1838 -136 1918 -132
rect 1838 -218 1842 -136
rect 1842 -218 1914 -136
rect 1914 -218 1918 -136
rect 1838 -222 1918 -218
rect -292 -826 -282 -762
rect -282 -826 -248 -762
rect -248 -826 -238 -762
rect 1684 -904 1782 -802
rect 1560 -988 1614 -982
rect 1560 -1032 1568 -988
rect 1568 -1032 1604 -988
rect 1604 -1032 1614 -988
rect 1560 -1034 1614 -1032
rect 2968 -942 3022 -940
rect 2968 -986 2978 -942
rect 2978 -986 3014 -942
rect 3014 -986 3022 -942
rect 2968 -1002 3022 -986
rect 764 -1238 820 -1236
rect 764 -1280 772 -1238
rect 772 -1280 810 -1238
rect 810 -1280 820 -1238
rect 764 -1290 820 -1280
rect 1838 -1234 1960 -1232
rect 1838 -1362 1842 -1234
rect 1842 -1362 1956 -1234
rect 1956 -1362 1960 -1234
rect 1838 -1366 1960 -1362
rect 914 -1682 966 -1506
rect 1432 -1680 1486 -1512
rect 2274 -1682 2328 -1494
rect 2792 -1684 2844 -1496
rect 522 -2418 574 -2414
rect 522 -2462 530 -2418
rect 530 -2462 566 -2418
rect 566 -2462 574 -2418
rect 522 -2466 574 -2462
rect 2828 -2418 2894 -2414
rect 2828 -2462 2832 -2418
rect 2832 -2462 2890 -2418
rect 2890 -2462 2894 -2418
rect 2828 -2466 2894 -2462
rect 1674 -2934 1726 -2882
rect 2368 -4294 2430 -4290
rect 2368 -4340 2374 -4294
rect 2374 -4340 2424 -4294
rect 2424 -4340 2430 -4294
rect 2368 -4344 2430 -4340
<< metal2 >>
rect -678 3068 -628 3244
rect -678 -404 -630 3068
rect 2162 2702 2248 2770
rect 2092 1722 2190 1728
rect 2092 1666 2108 1722
rect 2172 1666 2190 1722
rect 2092 1648 2190 1666
rect 2092 1576 3184 1648
rect 2974 204 3064 212
rect 692 198 3064 204
rect 692 190 1612 198
rect 692 -62 728 190
rect 784 -62 1612 190
rect 692 -66 1612 -62
rect 1664 -66 1744 198
rect 692 -70 1744 -66
rect 1800 196 2990 198
rect 1800 -66 2064 196
rect 2124 -66 2990 196
rect 1800 -70 2990 -66
rect 692 -72 2990 -70
rect 3044 -72 3064 198
rect 692 -76 3064 -72
rect 2974 -88 3064 -76
rect 94 -126 254 -120
rect 1800 -126 1960 -118
rect 94 -132 1960 -126
rect 94 -134 1838 -132
rect 94 -224 132 -134
rect 212 -222 1838 -134
rect 1918 -222 1960 -132
rect 212 -224 254 -222
rect 94 -232 254 -224
rect 1800 -230 1960 -222
rect -678 -452 1770 -404
rect 1722 -754 1770 -452
rect -298 -762 786 -756
rect -298 -826 -292 -762
rect -238 -826 786 -762
rect -298 -832 786 -826
rect 710 -1124 786 -832
rect 1678 -802 1788 -754
rect 1678 -904 1684 -802
rect 1782 -904 1788 -802
rect 1678 -920 1788 -904
rect 1964 -910 2074 -802
rect 2958 -940 3030 -936
rect 1544 -982 1628 -980
rect 1544 -1034 1560 -982
rect 1614 -1034 2162 -982
rect 1544 -1038 2162 -1034
rect 1544 -1040 1628 -1038
rect 710 -1200 1986 -1124
rect 1814 -1232 1986 -1200
rect 754 -1236 828 -1232
rect 754 -1290 764 -1236
rect 820 -1290 828 -1236
rect 754 -1300 828 -1290
rect 756 -2136 828 -1300
rect 1814 -1366 1838 -1232
rect 1960 -1366 1986 -1232
rect 1814 -1374 1986 -1366
rect 898 -1506 1500 -1490
rect 898 -1682 914 -1506
rect 966 -1512 1500 -1506
rect 966 -1680 1432 -1512
rect 1486 -1680 1500 -1512
rect 966 -1682 1500 -1680
rect 898 -1694 1500 -1682
rect 1460 -1696 1500 -1694
rect 514 -2208 828 -2136
rect 514 -2230 582 -2208
rect 512 -2410 582 -2230
rect 502 -2414 596 -2410
rect 502 -2466 522 -2414
rect 574 -2466 596 -2414
rect 502 -2470 596 -2466
rect 1658 -2878 1742 -2872
rect 1658 -2938 1670 -2878
rect 1730 -2938 1742 -2878
rect 1658 -2942 1742 -2938
rect 2106 -3032 2162 -1038
rect 2958 -1002 2968 -940
rect 3022 -1002 3030 -940
rect 3112 -1002 3184 1576
rect 2958 -1074 3184 -1002
rect 2260 -1494 2860 -1486
rect 2260 -1682 2274 -1494
rect 2328 -1496 2860 -1494
rect 2328 -1682 2792 -1496
rect 2260 -1684 2792 -1682
rect 2844 -1684 2860 -1496
rect 2260 -1690 2860 -1684
rect 2958 -2212 3030 -1074
rect 2866 -2278 3030 -2212
rect 2866 -2410 2932 -2278
rect 2798 -2414 2932 -2410
rect 2798 -2466 2828 -2414
rect 2894 -2466 2932 -2414
rect 2798 -2470 2932 -2466
rect 2106 -3088 2426 -3032
rect 2370 -4276 2426 -3088
rect 2360 -4290 2440 -4276
rect 2360 -4344 2368 -4290
rect 2430 -4344 2440 -4290
rect 2360 -4350 2440 -4344
rect 2378 -5478 2458 -5070
<< via2 >>
rect 1670 -2882 1730 -2878
rect 1670 -2934 1674 -2882
rect 1674 -2934 1726 -2882
rect 1726 -2934 1730 -2882
rect 1670 -2938 1730 -2934
<< metal3 >>
rect -704 3130 -604 3256
rect -1057 -922 2090 -796
rect -603 -5353 -477 -922
rect 1658 -2878 1742 -2872
rect 1658 -2938 1670 -2878
rect 1730 -2938 1742 -2878
rect 1658 -2942 1742 -2938
rect -603 -5479 3925 -5353
rect 3799 -7871 3925 -5479
<< metal4 >>
rect -704 3130 -604 3256
rect 1270 -3466 2134 -2118
rect 1316 -3472 1450 -3466
use sky130_fd_pr__cap_mim_m3_1_LABLLG  sky130_fd_pr__cap_mim_m3_1_LABLLG_0
timestamp 1702109072
transform 1 0 -17372 0 1 15572
box -16410 -15800 16410 15800
use sky130_fd_pr__cap_mim_m3_1_LABLLG  sky130_fd_pr__cap_mim_m3_1_LABLLG_1
timestamp 1702109072
transform 1 0 -17372 0 1 -16428
box -16410 -15800 16410 15800
use sky130_fd_pr__cap_mim_m3_1_S6JVQT  sky130_fd_pr__cap_mim_m3_1_S6JVQT_0
timestamp 1702106960
transform 0 -1 1670 1 0 -11886
box -6492 -2540 6492 2540
use sky130_fd_pr__cap_mim_m3_1_S6JVQT  sky130_fd_pr__cap_mim_m3_1_S6JVQT_1
timestamp 1702106960
transform 0 1 1670 -1 0 9178
box -6492 -2540 6492 2540
use sky130_fd_pr__cap_mim_m3_1_VYX8PH  sky130_fd_pr__cap_mim_m3_1_VYX8PH_0
timestamp 1702085311
transform 0 -1 1708 1 0 -3542
box -686 -540 686 540
use sky130_fd_pr__nfet_01v8_8BU2MY  sky130_fd_pr__nfet_01v8_8BU2MY_0
timestamp 1701653031
transform 1 0 1900 0 1 -1870
box -138 -226 138 226
use sky130_fd_pr__nfet_01v8_9GUA3Y  sky130_fd_pr__nfet_01v8_9GUA3Y_0
timestamp 1701652012
transform 1 0 504 0 1 -1470
box -138 -626 138 626
use sky130_fd_pr__nfet_01v8_9GUA3Y  sky130_fd_pr__nfet_01v8_9GUA3Y_1
timestamp 1701652012
transform 1 0 -156 0 1 -1470
box -138 -626 138 626
use sky130_fd_pr__nfet_01v8_HZDBC9  sky130_fd_pr__nfet_01v8_HZDBC9_0
timestamp 1701652675
transform 1 0 2559 0 1 -1470
box -287 -626 287 626
use sky130_fd_pr__nfet_01v8_HZDBC9  sky130_fd_pr__nfet_01v8_HZDBC9_1
timestamp 1701652675
transform 1 0 1201 0 1 -1470
box -287 -626 287 626
use sky130_fd_pr__pfet_01v8_AM3UTC  sky130_fd_pr__pfet_01v8_AM3UTC_0
timestamp 1701652012
transform 1 0 -156 0 1 260
box -174 -862 174 862
use sky130_fd_pr__pfet_01v8_AM3UTC  sky130_fd_pr__pfet_01v8_AM3UTC_1
timestamp 1701652012
transform 1 0 504 0 1 260
box -174 -862 174 862
use sky130_fd_pr__pfet_01v8_ESNC2G  sky130_fd_pr__pfet_01v8_ESNC2G_0
timestamp 1702085311
transform -1 0 2206 0 1 -2610
box -510 -162 510 162
use sky130_fd_pr__pfet_01v8_ESNC2G  sky130_fd_pr__pfet_01v8_ESNC2G_1
timestamp 1702085311
transform -1 0 3214 0 1 -2610
box -510 -162 510 162
use sky130_fd_pr__pfet_01v8_ESNC2G  sky130_fd_pr__pfet_01v8_ESNC2G_2
timestamp 1702085311
transform 1 0 186 0 1 -2610
box -510 -162 510 162
use sky130_fd_pr__pfet_01v8_ESNC2G  sky130_fd_pr__pfet_01v8_ESNC2G_3
timestamp 1702085311
transform 1 0 1194 0 1 -2610
box -510 -162 510 162
use sky130_fd_pr__pfet_01v8_ESNCXF  sky130_fd_pr__pfet_01v8_ESNCXF_0
timestamp 1702104985
transform 1 0 1090 0 1 -4494
box -460 -162 460 162
use sky130_fd_pr__pfet_01v8_ESNCXF  sky130_fd_pr__pfet_01v8_ESNCXF_1
timestamp 1702104985
transform -1 0 2090 0 1 -4494
box -460 -162 460 162
use sky130_fd_pr__pfet_01v8_ESNCXF  sky130_fd_pr__pfet_01v8_ESNCXF_2
timestamp 1702104985
transform -1 0 2090 0 1 -4934
box -460 -162 460 162
use sky130_fd_pr__pfet_01v8_ESNCXF  sky130_fd_pr__pfet_01v8_ESNCXF_3
timestamp 1702104985
transform 1 0 1090 0 1 -4934
box -460 -162 460 162
use sky130_fd_pr__pfet_01v8_ESNCXF  sky130_fd_pr__pfet_01v8_ESNCXF_4
timestamp 1702104985
transform 1 0 824 0 1 1866
box -460 -162 460 162
use sky130_fd_pr__pfet_01v8_ESNCXF  sky130_fd_pr__pfet_01v8_ESNCXF_5
timestamp 1702104985
transform -1 0 1824 0 1 1866
box -460 -162 460 162
use sky130_fd_pr__pfet_01v8_ESNCXF  sky130_fd_pr__pfet_01v8_ESNCXF_6
timestamp 1702104985
transform 1 0 824 0 1 2306
box -460 -162 460 162
use sky130_fd_pr__pfet_01v8_ESNCXF  sky130_fd_pr__pfet_01v8_ESNCXF_7
timestamp 1702104985
transform -1 0 1824 0 1 2306
box -460 -162 460 162
use sky130_fd_pr__pfet_01v8_S43UTC  sky130_fd_pr__pfet_01v8_S43UTC_0
timestamp 1701652012
transform 1 0 1880 0 1 660
box -174 -462 174 462
use sky130_fd_pr__pfet_01v8_S43UTC  sky130_fd_pr__pfet_01v8_S43UTC_1
timestamp 1701652012
transform 1 0 174 0 1 660
box -174 -462 174 462
use sky130_fd_pr__pfet_01v8_VBYK8W  sky130_fd_pr__pfet_01v8_VBYK8W_0
timestamp 1701652323
transform 1 0 1201 0 1 160
box -523 -962 523 962
use sky130_fd_pr__pfet_01v8_VBYK8W  sky130_fd_pr__pfet_01v8_VBYK8W_1
timestamp 1701652323
transform 1 0 2559 0 1 160
box -523 -962 523 962
<< labels >>
flabel viali -290 1206 -290 1206 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel via1 174 -182 174 -182 0 FreeSans 800 0 0 0 Vbias
port 4 nsew
flabel polycont 1730 -860 1730 -860 0 FreeSans 400 0 0 0 INP
port 5 nsew
flabel polycont 2020 -856 2020 -856 0 FreeSans 400 0 0 0 INN
port 6 nsew
flabel viali 1584 -1014 1584 -1014 0 FreeSans 400 0 0 0 V1N
port 7 nsew
flabel viali 3002 -970 3002 -970 0 FreeSans 400 0 0 0 V1P
port 8 nsew
flabel viali -164 -668 -164 -668 0 FreeSans 400 0 0 0 Vref
port 9 nsew
flabel polycont 500 -680 500 -680 0 FreeSans 400 0 0 0 Vcm_in
port 10 nsew
flabel viali -230 -2278 -230 -2278 0 FreeSans 800 0 0 0 VSS
port 11 nsew
flabel metal4 1638 -2622 1638 -2610 0 FreeSans 400 0 0 0 Vcm_out
port 12 nsew
<< end >>

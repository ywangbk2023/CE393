magic
tech sky130A
magscale 1 2
timestamp 1702063849
<< nwell >>
rect -410 1118 3356 1474
rect -410 1108 576 1118
rect 594 1108 638 1110
rect 658 1108 3356 1118
rect -410 1106 3356 1108
rect 594 1048 638 1106
rect 1972 1040 2006 1106
rect 42 264 88 272
rect 1748 268 1794 274
rect -40 134 -38 168
rect 10 104 342 264
rect 1746 204 1798 268
rect 1800 236 1960 254
rect 18 -524 330 104
rect 692 -76 3044 204
rect 1706 -80 2036 -76
rect 16 -602 346 -524
rect 470 -602 538 -524
rect 1724 -802 2036 -80
<< pmos >>
rect 470 -540 538 -524
<< ndiff >>
rect 1474 -1680 1486 -1666
rect 2274 -1604 2284 -1570
rect 2842 -1684 2844 -1496
<< poly >>
rect 94 -142 254 246
rect 94 -216 140 -142
rect 204 -216 254 -142
rect 94 -232 254 -216
rect 1800 -140 1960 254
rect 1800 -214 1846 -140
rect 1910 -214 1960 -140
rect 1800 -230 1960 -214
rect -184 -622 -136 -524
rect 470 -566 538 -540
rect 480 -622 528 -566
rect -194 -630 -126 -622
rect -194 -698 -178 -630
rect -142 -698 -126 -630
rect -194 -708 -126 -698
rect 470 -630 538 -622
rect 470 -698 486 -630
rect 522 -698 538 -630
rect 470 -708 538 -698
rect -76 -750 -8 -740
rect -124 -818 -60 -750
rect -24 -818 -8 -750
rect -124 -828 -8 -818
rect 356 -750 424 -740
rect 356 -818 372 -750
rect 408 -818 472 -750
rect 972 -756 1172 -708
rect 1230 -756 1430 -704
rect 356 -828 472 -818
rect 770 -762 1430 -756
rect 2330 -758 2530 -702
rect 2588 -758 2788 -696
rect 770 -818 1788 -762
rect 2330 -766 2788 -758
rect 770 -824 1694 -818
rect -124 -870 -76 -828
rect 424 -870 472 -828
rect 972 -830 1430 -824
rect 972 -870 1172 -830
rect 1230 -870 1430 -830
rect 1678 -894 1694 -824
rect 1772 -894 1788 -818
rect 1678 -910 1788 -894
rect 1964 -818 2990 -766
rect 1964 -894 1980 -818
rect 2058 -828 2990 -818
rect 2058 -894 2074 -828
rect 2330 -832 2788 -828
rect 2330 -862 2530 -832
rect 2588 -856 2788 -832
rect 1964 -910 2074 -894
rect 1820 -1240 1980 -1216
rect 1820 -1352 1848 -1240
rect 1948 -1352 1980 -1240
rect 1820 -1670 1980 -1352
<< polycont >>
rect 140 -216 204 -142
rect 1846 -214 1910 -140
rect -178 -698 -142 -630
rect 486 -698 522 -630
rect -60 -818 -24 -750
rect 372 -818 408 -750
rect 1694 -894 1772 -818
rect 1980 -894 2058 -818
rect 1848 -1352 1948 -1240
<< locali >>
rect 258 1352 308 1368
rect 258 1126 266 1352
rect 300 1126 308 1352
rect 258 1118 308 1126
rect 1960 1360 2022 1368
rect 1960 1124 1972 1360
rect 2006 1124 2022 1360
rect 1960 1118 2022 1124
rect 266 1042 300 1118
rect 1972 1040 2006 1118
rect -40 134 -38 168
rect 94 -138 254 -120
rect 94 -220 136 -138
rect 208 -220 254 -138
rect 94 -232 254 -220
rect 1800 -136 1960 -118
rect 1800 -218 1842 -136
rect 1914 -218 1960 -136
rect 1800 -230 1960 -218
rect -282 -756 -248 -544
rect -194 -630 -126 -622
rect -194 -698 -178 -630
rect -142 -698 -126 -630
rect -194 -708 -126 -698
rect 470 -630 538 -622
rect 470 -698 486 -630
rect 522 -698 538 -630
rect 470 -708 538 -698
rect -76 -750 -8 -740
rect 356 -750 424 -740
rect 596 -750 630 -544
rect -298 -762 -232 -756
rect -298 -826 -282 -762
rect -248 -826 -232 -762
rect -298 -832 -232 -826
rect -76 -818 -60 -750
rect -24 -818 372 -750
rect 408 -818 630 -750
rect -76 -828 -8 -818
rect 356 -828 424 -818
rect -282 -872 -248 -832
rect 596 -872 630 -818
rect 1184 -784 1218 -744
rect 1184 -826 1606 -784
rect 2542 -790 2576 -744
rect 1184 -876 1218 -826
rect 1184 -902 1218 -884
rect 1564 -982 1606 -826
rect 1678 -818 1788 -802
rect 1678 -894 1694 -818
rect 1772 -894 1788 -818
rect 1678 -910 1788 -894
rect 1964 -818 2074 -802
rect 1964 -894 1980 -818
rect 2058 -894 2074 -818
rect 2542 -832 3016 -790
rect 2542 -876 2576 -832
rect 1964 -910 2074 -894
rect 2974 -936 3016 -832
rect 2964 -942 3026 -936
rect 1554 -988 1616 -982
rect 1554 -1032 1568 -988
rect 1604 -1032 1616 -988
rect 2964 -986 2978 -942
rect 3014 -986 3026 -942
rect 2964 -992 3026 -986
rect 1554 -1038 1616 -1032
rect 1820 -1234 1980 -1216
rect 1820 -1362 1842 -1234
rect 1956 -1362 1980 -1234
rect 1820 -1374 1980 -1362
rect 2284 -1604 2286 -1570
rect 1774 -1868 1808 -1688
rect -64 -2118 -30 -2072
rect 378 -2118 412 -2072
rect 1992 -2118 2026 -1658
rect -72 -2124 -22 -2118
rect -72 -2360 -64 -2124
rect -30 -2360 -22 -2124
rect -72 -2368 -22 -2360
rect 370 -2124 420 -2118
rect 370 -2360 378 -2124
rect 412 -2360 420 -2124
rect 370 -2368 420 -2360
rect 1984 -2124 2034 -2118
rect 1984 -2360 1992 -2124
rect 2026 -2360 2034 -2124
rect 1984 -2368 2034 -2360
<< viali >>
rect 266 1126 300 1352
rect 1972 1124 2006 1360
rect 136 -142 208 -138
rect 136 -216 140 -142
rect 140 -216 204 -142
rect 204 -216 208 -142
rect 136 -220 208 -216
rect 1842 -140 1914 -136
rect 1842 -214 1846 -140
rect 1846 -214 1910 -140
rect 1910 -214 1914 -140
rect 1842 -218 1914 -214
rect -178 -682 -142 -648
rect -282 -826 -248 -762
rect 1568 -1032 1604 -988
rect 2978 -986 3014 -942
rect 1842 -1240 1956 -1234
rect 1842 -1352 1848 -1240
rect 1848 -1352 1948 -1240
rect 1948 -1352 1956 -1240
rect 1842 -1362 1956 -1352
rect -64 -2360 -30 -2124
rect 378 -2360 412 -2124
rect 1992 -2360 2026 -2124
<< metal1 >>
rect -346 1360 3250 1368
rect -346 1352 1972 1360
rect -346 1126 266 1352
rect 300 1126 1972 1352
rect -346 1124 1972 1126
rect 2006 1124 3250 1360
rect -346 1118 3250 1124
rect 42 216 88 272
rect -30 118 384 216
rect 1748 204 1794 274
rect 714 190 808 204
rect 714 -62 728 190
rect 784 -62 808 190
rect 714 -76 808 -62
rect 1590 198 1682 204
rect 1590 -66 1612 198
rect 1664 -66 1682 198
rect 1590 -76 1682 -66
rect 1732 198 1808 204
rect 1732 -70 1744 198
rect 1800 -70 1808 198
rect 1732 -76 1808 -70
rect 2056 196 2084 204
rect 2974 198 3064 212
rect 2056 -66 2064 196
rect 2056 -76 2084 -66
rect 2974 -72 2990 198
rect 3044 -72 3064 198
rect 2974 -88 3064 -72
rect 94 -134 254 -120
rect 94 -224 132 -134
rect 212 -224 254 -134
rect 94 -232 254 -224
rect 1800 -132 1960 -118
rect 1800 -222 1838 -132
rect 1918 -222 1960 -132
rect 1800 -230 1960 -222
rect -296 -648 -116 -642
rect -296 -682 -178 -648
rect -142 -682 -116 -648
rect -296 -690 -116 -682
rect -298 -762 -232 -756
rect -298 -826 -292 -762
rect -238 -826 -232 -762
rect -298 -832 -232 -826
rect 2954 -942 3038 -936
rect 1544 -988 1628 -982
rect 1544 -1032 1568 -988
rect 1604 -1032 1628 -988
rect 2954 -986 2978 -942
rect 3014 -986 3038 -942
rect 2954 -992 3038 -986
rect 1544 -1038 1628 -1032
rect 1814 -1232 1986 -1216
rect 1814 -1366 1838 -1232
rect 1960 -1366 1986 -1232
rect 1814 -1374 1986 -1366
rect 1652 -1486 2322 -1450
rect 906 -1506 984 -1490
rect 906 -1682 914 -1506
rect 966 -1682 984 -1506
rect 906 -1694 984 -1682
rect 1418 -1512 1500 -1490
rect 1418 -1680 1432 -1512
rect 1486 -1680 1500 -1512
rect 1418 -1694 1500 -1680
rect 1460 -1696 1500 -1694
rect 1652 -1494 2336 -1486
rect 1652 -1612 2274 -1494
rect 1652 -1730 1814 -1612
rect 2268 -1682 2274 -1612
rect 2328 -1682 2336 -1494
rect 2268 -1690 2336 -1682
rect 2788 -1496 2860 -1486
rect 2788 -1684 2792 -1496
rect 2844 -1684 2860 -1496
rect 2788 -1690 2860 -1684
rect 1472 -1882 1814 -1730
rect -326 -2124 3294 -2118
rect -326 -2360 -64 -2124
rect -30 -2360 378 -2124
rect 412 -2360 1992 -2124
rect 2026 -2360 3294 -2124
rect -326 -2368 3294 -2360
<< via1 >>
rect 728 -62 784 190
rect 1612 -66 1664 198
rect 1744 -70 1800 198
rect 2064 -66 2124 196
rect 2990 -72 3044 198
rect 132 -138 212 -134
rect 132 -220 136 -138
rect 136 -220 208 -138
rect 208 -220 212 -138
rect 132 -224 212 -220
rect 1838 -136 1918 -132
rect 1838 -218 1842 -136
rect 1842 -218 1914 -136
rect 1914 -218 1918 -136
rect 1838 -222 1918 -218
rect -292 -826 -282 -762
rect -282 -826 -248 -762
rect -248 -826 -238 -762
rect 1838 -1234 1960 -1232
rect 1838 -1362 1842 -1234
rect 1842 -1362 1956 -1234
rect 1956 -1362 1960 -1234
rect 1838 -1366 1960 -1362
rect 914 -1682 966 -1506
rect 1432 -1680 1486 -1512
rect 2274 -1682 2328 -1494
rect 2792 -1684 2844 -1496
<< metal2 >>
rect 2974 204 3064 212
rect 692 198 3064 204
rect 692 190 1612 198
rect 692 -62 728 190
rect 784 -62 1612 190
rect 692 -66 1612 -62
rect 1664 -66 1744 198
rect 692 -70 1744 -66
rect 1800 196 2990 198
rect 1800 -66 2064 196
rect 2124 -66 2990 196
rect 1800 -70 2990 -66
rect 692 -72 2990 -70
rect 3044 -72 3064 198
rect 692 -76 3064 -72
rect 2974 -88 3064 -76
rect 94 -126 254 -120
rect 1800 -126 1960 -118
rect 94 -132 1960 -126
rect 94 -134 1838 -132
rect 94 -224 132 -134
rect 212 -222 1838 -134
rect 1918 -222 1960 -132
rect 212 -224 254 -222
rect 94 -232 254 -224
rect 1800 -230 1960 -222
rect -298 -762 786 -756
rect -298 -826 -292 -762
rect -238 -826 786 -762
rect -298 -832 786 -826
rect 710 -1124 786 -832
rect 710 -1200 1986 -1124
rect 1814 -1232 1986 -1200
rect 1814 -1366 1838 -1232
rect 1960 -1366 1986 -1232
rect 1814 -1374 1986 -1366
rect 898 -1506 1500 -1490
rect 898 -1682 914 -1506
rect 966 -1512 1500 -1506
rect 966 -1680 1432 -1512
rect 1486 -1680 1500 -1512
rect 966 -1682 1500 -1680
rect 898 -1694 1500 -1682
rect 2260 -1494 2860 -1486
rect 2260 -1682 2274 -1494
rect 2328 -1496 2860 -1494
rect 2328 -1682 2792 -1496
rect 2260 -1684 2792 -1682
rect 2844 -1684 2860 -1496
rect 2260 -1690 2860 -1684
rect 1460 -1696 1500 -1694
use sky130_fd_pr__nfet_01v8_8BU2MY  sky130_fd_pr__nfet_01v8_8BU2MY_0
timestamp 1701653031
transform 1 0 1900 0 1 -1870
box -138 -226 138 226
use sky130_fd_pr__nfet_01v8_9GUA3Y  sky130_fd_pr__nfet_01v8_9GUA3Y_0
timestamp 1701652012
transform 1 0 504 0 1 -1470
box -138 -626 138 626
use sky130_fd_pr__nfet_01v8_9GUA3Y  sky130_fd_pr__nfet_01v8_9GUA3Y_1
timestamp 1701652012
transform 1 0 -156 0 1 -1470
box -138 -626 138 626
use sky130_fd_pr__nfet_01v8_HZDBC9  sky130_fd_pr__nfet_01v8_HZDBC9_0
timestamp 1701652675
transform 1 0 2559 0 1 -1470
box -287 -626 287 626
use sky130_fd_pr__nfet_01v8_HZDBC9  sky130_fd_pr__nfet_01v8_HZDBC9_1
timestamp 1701652675
transform 1 0 1201 0 1 -1470
box -287 -626 287 626
use sky130_fd_pr__pfet_01v8_AM3UTC  sky130_fd_pr__pfet_01v8_AM3UTC_0
timestamp 1701652012
transform 1 0 -156 0 1 260
box -174 -862 174 862
use sky130_fd_pr__pfet_01v8_AM3UTC  sky130_fd_pr__pfet_01v8_AM3UTC_1
timestamp 1701652012
transform 1 0 504 0 1 260
box -174 -862 174 862
use sky130_fd_pr__pfet_01v8_S43UTC  sky130_fd_pr__pfet_01v8_S43UTC_0
timestamp 1701652012
transform 1 0 1880 0 1 660
box -174 -462 174 462
use sky130_fd_pr__pfet_01v8_S43UTC  sky130_fd_pr__pfet_01v8_S43UTC_1
timestamp 1701652012
transform 1 0 174 0 1 660
box -174 -462 174 462
use sky130_fd_pr__pfet_01v8_VBYK8W  sky130_fd_pr__pfet_01v8_VBYK8W_0
timestamp 1701652323
transform 1 0 1201 0 1 160
box -523 -962 523 962
use sky130_fd_pr__pfet_01v8_VBYK8W  sky130_fd_pr__pfet_01v8_VBYK8W_1
timestamp 1701652323
transform 1 0 2559 0 1 160
box -523 -962 523 962
<< end >>

magic
tech sky130A
timestamp 1702099645
<< nwell >>
rect 424 247 525 248
<< nmos >>
rect 300 41 324 141
rect 353 41 377 141
rect 571 -59 595 141
rect 624 -59 648 141
rect 733 -59 757 141
<< ndiff >>
rect 271 135 300 141
rect 271 47 277 135
rect 294 47 300 135
rect 271 41 300 47
rect 324 135 353 141
rect 324 47 330 135
rect 347 47 353 135
rect 324 41 353 47
rect 377 135 406 141
rect 377 47 383 135
rect 400 47 406 135
rect 377 41 406 47
rect 542 135 571 141
rect 542 -53 548 135
rect 565 -53 571 135
rect 542 -59 571 -53
rect 595 135 624 141
rect 595 -53 601 135
rect 618 -53 624 135
rect 595 -59 624 -53
rect 648 135 677 141
rect 648 -53 654 135
rect 671 -53 677 135
rect 648 -59 677 -53
rect 704 135 733 141
rect 704 -53 710 135
rect 727 -53 733 135
rect 704 -59 733 -53
rect 757 135 786 141
rect 757 -53 763 135
rect 780 -53 786 135
rect 757 -59 786 -53
<< ndiffc >>
rect 277 47 294 135
rect 330 47 347 135
rect 383 47 400 135
rect 548 -53 565 135
rect 601 -53 618 135
rect 654 -53 671 135
rect 710 -53 727 135
rect 763 -53 780 135
<< poly >>
rect -472 515 -421 523
rect -472 479 -464 515
rect -430 479 -421 515
rect -472 472 -421 479
rect -471 440 -446 472
rect 138 153 163 266
rect 191 152 215 276
rect 300 141 324 273
rect 353 141 377 273
rect 462 149 486 273
rect 571 141 595 273
rect 624 141 648 273
rect 733 141 757 267
rect 137 18 162 28
rect 105 9 162 18
rect 105 -16 115 9
rect 138 -15 162 9
rect 191 22 215 28
rect 300 22 324 41
rect 191 15 239 22
rect 191 -6 212 15
rect 231 -6 239 15
rect 191 -13 239 -6
rect 289 16 324 22
rect 289 -1 298 16
rect 316 -1 324 16
rect 289 -9 324 -1
rect 353 21 377 41
rect 462 29 479 31
rect 353 14 388 21
rect 353 -3 361 14
rect 380 -3 388 14
rect 353 -10 388 -3
rect 456 -1 491 29
rect 138 -16 147 -15
rect 105 -24 147 -16
rect 456 -18 464 -1
rect 483 -18 491 -1
rect 456 -26 491 -18
rect 571 -71 595 -59
rect 624 -71 648 -59
rect 733 -71 757 -59
rect 565 -98 600 -71
rect 565 -115 573 -98
rect 592 -115 600 -98
rect 565 -123 600 -115
rect 624 -101 659 -71
rect 624 -118 632 -101
rect 651 -118 659 -101
rect 624 -125 659 -118
rect 733 -100 768 -71
rect 733 -117 741 -100
rect 760 -117 768 -100
rect 733 -124 768 -117
<< polycont >>
rect -464 479 -430 515
rect 115 -16 138 9
rect 212 -6 231 15
rect 298 -1 316 16
rect 361 -3 380 14
rect 464 -18 483 -1
rect 573 -115 592 -98
rect 632 -118 651 -101
rect 741 -117 760 -100
<< locali >>
rect 6356 1489 6428 1497
rect 6356 1435 6364 1489
rect 6420 1435 6428 1489
rect 6356 1428 6428 1435
rect -472 515 -421 523
rect -472 479 -464 515
rect -430 479 -421 515
rect -472 472 -421 479
rect 548 472 565 509
rect 654 472 671 481
rect 763 475 780 492
rect 115 380 132 381
rect 221 380 238 381
rect 277 380 294 382
rect 383 379 400 382
rect 492 381 509 387
rect -251 298 -208 304
rect -251 272 -241 298
rect -216 272 -208 298
rect -251 266 -208 272
rect -318 240 -276 246
rect -244 240 -213 266
rect 168 241 185 276
rect 330 241 347 277
rect 439 241 456 277
rect 601 241 618 276
rect 710 241 727 276
rect 90 240 804 241
rect -440 237 804 240
rect -440 236 -311 237
rect -441 219 -311 236
rect -318 207 -311 219
rect -283 222 804 237
rect -283 219 93 222
rect -283 207 -276 219
rect -318 199 -276 207
rect -65 167 804 187
rect -65 166 115 167
rect 168 143 185 167
rect 277 135 294 143
rect 277 39 294 47
rect 330 135 347 167
rect 439 143 456 167
rect 330 39 347 47
rect 383 135 400 143
rect 383 39 400 47
rect 548 135 565 143
rect 115 38 132 39
rect 492 38 509 39
rect 105 9 147 18
rect 105 -16 115 9
rect 138 -16 147 9
rect 204 15 239 22
rect 204 -6 212 15
rect 231 -6 239 15
rect 204 -13 239 -6
rect 289 16 324 22
rect 289 -1 298 16
rect 316 -1 324 16
rect 289 -9 324 -1
rect 353 14 388 21
rect 353 -3 361 14
rect 380 -3 388 14
rect 353 -10 388 -3
rect 456 -1 491 6
rect 105 -24 147 -16
rect 456 -18 464 -1
rect 483 -18 491 -1
rect 456 -26 491 -18
rect 548 -61 565 -53
rect 601 135 618 167
rect 601 -61 618 -53
rect 654 135 671 143
rect 654 -63 671 -53
rect 710 135 727 167
rect 710 -63 727 -53
rect 763 135 780 143
rect 763 -64 780 -53
rect 565 -98 600 -91
rect 565 -115 573 -98
rect 592 -115 600 -98
rect 565 -123 600 -115
rect 624 -101 659 -93
rect 624 -118 632 -101
rect 651 -118 659 -101
rect 624 -125 659 -118
rect 733 -100 768 -92
rect 733 -117 741 -100
rect 760 -117 768 -100
rect 733 -124 768 -117
<< viali >>
rect 6364 1435 6420 1489
rect -241 272 -216 298
rect -311 207 -283 237
rect 277 47 294 135
rect 330 47 347 135
rect 383 47 400 135
rect 548 -53 565 135
rect 601 -53 618 135
rect 654 -53 671 135
rect 710 -53 727 135
rect 763 -53 780 135
<< metal1 >>
rect 6356 1489 6429 1501
rect -3296 1453 -3250 1458
rect -3296 1416 -3291 1453
rect -3255 1416 -3250 1453
rect 6356 1435 6364 1489
rect 6420 1435 6429 1489
rect 6356 1428 6429 1435
rect -3296 1376 -3250 1416
rect -3403 1059 -3350 1136
rect -3403 1024 -3395 1059
rect -3358 1024 -3350 1059
rect -3403 390 -3350 1024
rect -3295 965 -3253 1376
rect -915 1087 -863 1094
rect -1688 1058 -1613 1069
rect -1688 1004 -1678 1058
rect -1624 1004 -1613 1058
rect -915 1053 -907 1087
rect -870 1053 -863 1087
rect -542 1079 -490 1086
rect -542 1075 -536 1079
rect -915 1047 -863 1053
rect -1688 994 -1613 1004
rect -3295 541 -3250 965
rect -1678 668 -1614 994
rect -908 741 -871 1047
rect -544 1042 -536 1075
rect -497 1042 -490 1079
rect -544 1037 -490 1042
rect -544 807 -495 1037
rect -101 907 -54 910
rect -101 883 -47 907
rect -101 847 -96 883
rect -59 861 -47 883
rect -59 847 -44 861
rect -101 843 -44 847
rect -544 794 -132 807
rect -544 772 -128 794
rect -537 769 -128 772
rect -908 738 -203 741
rect -908 697 -200 738
rect -887 696 -855 697
rect -310 668 -279 672
rect -1698 625 -279 668
rect -499 541 -474 542
rect -3295 487 -474 541
rect -3295 480 -3250 487
rect -2621 390 -729 393
rect -3403 336 -729 390
rect -499 383 -474 487
rect -310 400 -279 625
rect -240 447 -200 697
rect -168 497 -128 769
rect -84 545 -44 843
rect 707 567 754 577
rect 707 551 714 567
rect -85 543 39 545
rect -85 516 402 543
rect -85 513 39 516
rect -168 493 -27 497
rect -168 466 296 493
rect -168 465 -27 466
rect -168 464 -59 465
rect -240 445 -130 447
rect -240 418 238 445
rect -240 417 -130 418
rect -239 415 -130 417
rect 114 401 134 403
rect -249 400 134 401
rect -310 374 134 400
rect -310 372 -210 374
rect 114 338 134 374
rect 221 371 238 418
rect 276 341 296 466
rect 382 338 402 516
rect 544 532 714 551
rect 748 551 754 567
rect 748 532 757 551
rect 544 520 757 532
rect 544 518 732 520
rect 544 505 571 518
rect 543 501 571 505
rect 733 501 791 502
rect 543 460 570 501
rect 651 500 1676 501
rect 650 475 1676 500
rect 467 454 512 460
rect 650 455 677 475
rect 467 419 474 454
rect 506 419 512 454
rect 467 406 512 419
rect 489 375 512 406
rect 1630 447 1676 475
rect 1630 411 1635 447
rect 1670 411 1676 447
rect 1630 405 1676 411
rect 3260 467 3319 474
rect 3260 430 3270 467
rect 3308 430 3319 467
rect -3403 333 -1511 336
rect -786 164 -732 336
rect -251 298 -207 304
rect -251 272 -241 298
rect -216 272 -207 298
rect -251 266 -207 272
rect -318 237 -275 245
rect -318 207 -311 237
rect -283 207 -275 237
rect -318 164 -275 207
rect 115 203 132 314
rect 114 176 133 203
rect -786 121 -275 164
rect -318 114 -275 121
rect 115 110 132 176
rect 221 112 238 316
rect 277 141 294 324
rect 383 141 400 324
rect 274 135 297 141
rect 274 47 277 135
rect 294 47 297 135
rect 274 41 297 47
rect 327 135 350 141
rect 327 47 330 135
rect 347 47 350 135
rect 327 41 350 47
rect 380 135 403 141
rect 380 47 383 135
rect 400 47 403 135
rect 492 118 509 322
rect 548 141 565 318
rect 654 141 671 317
rect 763 238 780 314
rect 3260 238 3319 430
rect 763 193 3319 238
rect 763 141 780 193
rect 545 135 568 141
rect 380 41 403 47
rect 545 -53 548 135
rect 565 -53 568 135
rect 545 -59 568 -53
rect 598 135 621 141
rect 598 -53 601 135
rect 618 -53 621 135
rect 598 -59 621 -53
rect 651 135 674 141
rect 651 -53 654 135
rect 671 -53 674 135
rect 651 -59 674 -53
rect 707 135 730 141
rect 707 -53 710 135
rect 727 -53 730 135
rect 707 -59 730 -53
rect 760 135 783 141
rect 760 -53 763 135
rect 780 -53 783 135
rect 760 -59 783 -53
<< via1 >>
rect -3291 1416 -3255 1453
rect 6364 1436 6420 1489
rect -3395 1024 -3358 1059
rect -1678 1004 -1624 1058
rect -907 1053 -870 1087
rect -536 1042 -497 1079
rect -96 847 -59 883
rect 714 532 748 567
rect 474 419 506 454
rect 1635 411 1670 447
rect 3270 430 3308 467
<< metal2 >>
rect 6357 1489 6428 1498
rect -3296 1453 -3249 1458
rect -3296 1415 -3291 1453
rect -3255 1415 -3249 1453
rect 6357 1435 6364 1489
rect 6420 1435 6428 1489
rect 6357 1430 6428 1435
rect -3296 1410 -3249 1415
rect -915 1087 -863 1094
rect -3402 1059 -3350 1068
rect -3402 1024 -3395 1059
rect -3358 1024 -3350 1059
rect -3402 1018 -3350 1024
rect -1688 1059 -1613 1069
rect -1688 1002 -1679 1059
rect -1624 1002 -1613 1059
rect -915 1052 -907 1087
rect -870 1052 -863 1087
rect -915 1047 -863 1052
rect -542 1079 -490 1086
rect -542 1042 -536 1079
rect -497 1042 -490 1079
rect -542 1037 -490 1042
rect -1688 994 -1613 1002
rect -101 883 -54 889
rect -101 847 -97 883
rect -59 847 -54 883
rect -101 842 -54 847
rect 706 567 756 577
rect 706 566 714 567
rect 706 532 713 566
rect 748 537 756 567
rect 748 532 755 537
rect 706 524 755 532
rect 3260 467 3316 474
rect 467 454 512 460
rect 467 419 474 454
rect 506 419 512 454
rect 467 413 512 419
rect 1630 447 1676 454
rect 1630 411 1634 447
rect 1670 411 1676 447
rect 3260 430 3270 467
rect 3308 430 3316 467
rect 3260 423 3316 430
rect 1630 405 1676 411
<< via2 >>
rect -3291 1416 -3255 1453
rect -3291 1415 -3255 1416
rect 6364 1436 6420 1489
rect 6364 1435 6420 1436
rect -3395 1024 -3358 1059
rect -1679 1058 -1624 1059
rect -1679 1004 -1678 1058
rect -1678 1004 -1624 1058
rect -1679 1002 -1624 1004
rect -907 1053 -870 1087
rect -907 1052 -870 1053
rect -536 1042 -497 1079
rect -97 847 -96 883
rect -96 847 -59 883
rect 713 532 714 566
rect 714 532 748 566
rect 474 419 506 454
rect 1634 411 1635 447
rect 1635 411 1670 447
rect 3270 430 3308 467
<< metal3 >>
rect -3691 1496 -3154 1503
rect 5848 1496 6427 1497
rect -3691 1489 6427 1496
rect -3691 1453 6364 1489
rect -3691 1415 -3291 1453
rect -3255 1435 6364 1453
rect 6420 1435 6427 1489
rect -3255 1431 6427 1435
rect -3255 1415 -3134 1431
rect -3691 1411 -3134 1415
rect -3690 1255 -3651 1411
rect -3296 1410 -3249 1411
rect -3173 1246 -3134 1411
rect -2754 1249 -2715 1330
rect -2383 1248 -2344 1334
rect -1964 1253 -1925 1340
rect -1585 1255 -1546 1431
rect -1200 1261 -1161 1344
rect -823 1257 -784 1431
rect -403 1264 -364 1431
rect 34 1277 73 1431
rect 480 1266 519 1431
rect 880 1275 919 1431
rect 1330 1281 1369 1431
rect 1718 1281 1757 1431
rect 2111 1288 2150 1431
rect 2503 1292 2542 1431
rect 2958 1283 2997 1431
rect 3354 1279 3393 1431
rect 3747 1281 3786 1431
rect 4146 1281 4185 1431
rect 4537 1281 4576 1431
rect 4925 1283 4964 1431
rect 5325 1281 5364 1431
rect 5717 1287 5756 1431
rect 5848 1430 6427 1431
rect 6356 1429 6427 1430
rect -2873 1147 -2712 1178
rect -2456 1149 -2295 1180
rect -2074 1150 -1913 1181
rect -3402 1059 -3350 1137
rect -1682 1069 -1627 1158
rect -1290 1153 -1129 1184
rect -915 1123 -864 1129
rect -915 1087 -862 1123
rect -3402 1024 -3395 1059
rect -3358 1024 -3350 1059
rect -3402 1018 -3350 1024
rect -1688 1059 -1613 1069
rect -1688 1001 -1679 1059
rect -1624 1001 -1613 1059
rect -915 1052 -907 1087
rect -870 1076 -862 1087
rect -542 1080 -490 1147
rect -870 1052 -863 1076
rect -915 1047 -863 1052
rect -542 1042 -536 1080
rect -497 1042 -490 1080
rect -542 1037 -490 1042
rect -1688 994 -1613 1001
rect -101 883 -54 943
rect -101 847 -97 883
rect -59 847 -54 883
rect -101 842 -54 847
rect 705 567 758 577
rect 346 460 389 566
rect 705 532 713 567
rect 748 532 758 567
rect 705 521 758 532
rect 3260 467 3316 474
rect 346 454 524 460
rect 346 419 474 454
rect 506 419 524 454
rect 346 412 524 419
rect 1626 447 1680 457
rect 1626 411 1633 447
rect 1671 411 1680 447
rect 3260 430 3270 467
rect 3308 430 3316 467
rect 3260 423 3316 430
rect 1626 399 1680 411
<< via3 >>
rect -3291 1415 -3255 1453
rect 6364 1435 6420 1489
rect -3395 1024 -3358 1059
rect -1679 1002 -1624 1059
rect -1679 1001 -1624 1002
rect -907 1052 -870 1087
rect -536 1079 -497 1080
rect -536 1042 -497 1079
rect -97 847 -59 883
rect 713 566 748 567
rect 713 532 748 566
rect 474 419 506 454
rect 1633 411 1634 447
rect 1634 411 1670 447
rect 1670 411 1671 447
rect 3270 430 3308 467
<< metal4 >>
rect -3691 1496 -3154 1503
rect 5848 1496 6427 1497
rect -3691 1489 6427 1496
rect -3691 1453 6364 1489
rect -3691 1415 -3291 1453
rect -3255 1435 6364 1453
rect 6420 1435 6427 1489
rect -3255 1431 6427 1435
rect -3255 1415 -3134 1431
rect -3691 1411 -3134 1415
rect -3690 1255 -3651 1411
rect -3173 1246 -3134 1411
rect -2754 1249 -2715 1330
rect -2383 1248 -2344 1334
rect -1964 1253 -1925 1340
rect -1585 1255 -1546 1431
rect -1200 1261 -1161 1344
rect -823 1257 -784 1431
rect -403 1264 -364 1431
rect 34 1277 73 1431
rect 480 1266 519 1431
rect 880 1275 919 1431
rect 1330 1281 1369 1431
rect 1718 1281 1757 1431
rect 2111 1288 2150 1431
rect 2503 1292 2542 1431
rect 2958 1283 2997 1431
rect 3354 1279 3393 1431
rect 3747 1281 3786 1431
rect 4146 1281 4185 1431
rect 4537 1281 4576 1431
rect 4925 1283 4964 1431
rect 5325 1281 5364 1431
rect 5717 1287 5756 1431
rect 5848 1430 6427 1431
rect -2873 1147 -2712 1178
rect -2456 1149 -2295 1180
rect -2074 1150 -1913 1181
rect -3402 1059 -3350 1137
rect -1682 1069 -1627 1158
rect -1290 1153 -1129 1184
rect -915 1123 -864 1129
rect -915 1087 -862 1123
rect -3402 1024 -3395 1059
rect -3358 1024 -3350 1059
rect -3402 1018 -3350 1024
rect -1688 1059 -1613 1069
rect -1688 1001 -1679 1059
rect -1624 1001 -1613 1059
rect -915 1052 -907 1087
rect -870 1076 -862 1087
rect -542 1080 -490 1147
rect -870 1052 -864 1076
rect -915 1047 -864 1052
rect -542 1042 -536 1080
rect -497 1042 -490 1080
rect -542 1037 -490 1042
rect -1688 994 -1613 1001
rect -101 883 -54 943
rect -101 847 -97 883
rect -59 847 -54 883
rect -101 843 -54 847
rect 706 576 755 577
rect 705 567 757 576
rect 346 460 389 566
rect 705 532 713 567
rect 748 532 757 567
rect 705 521 757 532
rect 346 454 524 460
rect 346 419 474 454
rect 506 419 524 454
rect 708 459 756 521
rect 788 459 836 598
rect 1182 547 1230 596
rect 1182 546 1231 547
rect 1183 467 1231 546
rect 1635 501 1676 605
rect 1183 459 1233 467
rect 708 419 1233 459
rect 346 412 524 419
rect 732 417 1233 419
rect 1631 454 1676 501
rect 2029 454 2070 610
rect 2424 454 2465 608
rect 2820 454 2861 605
rect 3266 474 3307 606
rect 3661 474 3702 610
rect 4056 474 4097 622
rect 4451 474 4492 618
rect 4846 474 4887 613
rect 5242 474 5283 601
rect 5637 474 5678 610
rect 6031 474 6072 606
rect 3265 467 6072 474
rect 1631 447 2864 454
rect 1631 411 1633 447
rect 1671 411 2864 447
rect 3265 430 3270 467
rect 3308 430 6072 467
rect 3265 426 6072 430
rect 1631 407 2864 411
rect 1631 406 1676 407
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_0
timestamp 1701930086
transform 1 0 191 0 1 950
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_1
timestamp 1701930086
transform 1 0 637 0 1 950
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_2
timestamp 1701930086
transform 1 0 1032 0 1 950
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_3
timestamp 1701930086
transform 1 0 5875 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_4
timestamp 1701930086
transform 1 0 4690 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_5
timestamp 1701930086
transform 1 0 5085 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_6
timestamp 1701930086
transform 1 0 5480 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_7
timestamp 1701930086
transform 1 0 2268 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_8
timestamp 1701930086
transform 1 0 2663 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_9
timestamp 1701930086
transform 1 0 1873 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_10
timestamp 1701930086
transform 1 0 1478 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_11
timestamp 1701930086
transform 1 0 3109 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_12
timestamp 1701930086
transform 1 0 3504 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_13
timestamp 1701930086
transform 1 0 4294 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_7AZ2EY  sky130_fd_pr__cap_mim_m3_1_7AZ2EY_14
timestamp 1701930086
transform 1 0 3899 0 1 957
box -203 -420 203 420
use sky130_fd_pr__cap_mim_m3_1_76Y692  sky130_fd_pr__cap_mim_m3_1_76Y692_0
timestamp 1701930086
transform 1 0 -250 0 1 1145
box -198 -220 198 220
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_0
timestamp 1701930086
transform 1 0 -1817 0 1 1227
box -193 -120 193 120
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_1
timestamp 1701930086
transform 1 0 -2608 0 1 1225
box -193 -120 193 120
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_2
timestamp 1701930086
transform 1 0 -3024 0 1 1224
box -193 -120 193 120
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_3
timestamp 1701930086
transform 1 0 -3540 0 1 1223
box -193 -120 193 120
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_4
timestamp 1701930086
transform 1 0 -1442 0 1 1228
box -193 -120 193 120
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_5
timestamp 1701930086
transform 1 0 -2233 0 1 1226
box -193 -120 193 120
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_6
timestamp 1701930086
transform 1 0 -1056 0 1 1226
box -193 -120 193 120
use sky130_fd_pr__cap_mim_m3_1_FJFAMD  sky130_fd_pr__cap_mim_m3_1_FJFAMD_7
timestamp 1701930086
transform 1 0 -681 0 1 1227
box -193 -120 193 120
use sky130_fd_pr__nfet_01v8_NQT7YS  sky130_fd_pr__nfet_01v8_NQT7YS_0
timestamp 1701909091
transform 1 0 474 0 1 91
box -41 -63 41 63
use sky130_fd_pr__nfet_01v8_NQT7YS  sky130_fd_pr__nfet_01v8_NQT7YS_1
timestamp 1701909091
transform 1 0 150 0 1 91
box -41 -63 41 63
use sky130_fd_pr__nfet_01v8_NQT7YS  sky130_fd_pr__nfet_01v8_NQT7YS_2
timestamp 1701909091
transform 1 0 203 0 1 91
box -41 -63 41 63
use sky130_fd_pr__pfet_01v8_A7S2BQ  sky130_fd_pr__pfet_01v8_A7S2BQ_0
timestamp 1702062038
transform 1 0 -459 0 1 328
box -59 -131 59 131
use sky130_fd_pr__pfet_01v8_A7S2BQ  sky130_fd_pr__pfet_01v8_A7S2BQ_1
timestamp 1702062038
transform 1 0 636 0 1 378
box -59 -131 59 131
use sky130_fd_pr__pfet_01v8_A7S2BQ  sky130_fd_pr__pfet_01v8_A7S2BQ_2
timestamp 1702062038
transform 1 0 583 0 1 378
box -59 -131 59 131
use sky130_fd_pr__pfet_01v8_A7S2BQ  sky130_fd_pr__pfet_01v8_A7S2BQ_3
timestamp 1702062038
transform 1 0 745 0 1 378
box -59 -131 59 131
use sky130_fd_pr__pfet_01v8_AZSHBQ  sky130_fd_pr__pfet_01v8_AZSHBQ_0
timestamp 1701909091
transform 1 0 312 0 1 328
box -59 -81 59 81
use sky130_fd_pr__pfet_01v8_AZSHBQ  sky130_fd_pr__pfet_01v8_AZSHBQ_1
timestamp 1701909091
transform 1 0 365 0 1 328
box -59 -81 59 81
use sky130_fd_pr__pfet_01v8_AZSHBQ  sky130_fd_pr__pfet_01v8_AZSHBQ_2
timestamp 1701909091
transform 1 0 150 0 1 328
box -59 -81 59 81
use sky130_fd_pr__pfet_01v8_AZSHBQ  sky130_fd_pr__pfet_01v8_AZSHBQ_3
timestamp 1701909091
transform 1 0 203 0 1 328
box -59 -81 59 81
use sky130_fd_pr__pfet_01v8_AZSHBQ  sky130_fd_pr__pfet_01v8_AZSHBQ_4
timestamp 1701909091
transform 1 0 474 0 1 329
box -59 -81 59 81
<< labels >>
flabel poly 733 -123 768 -91 0 FreeSans 8 0 0 0 Sw7
flabel space 844 -74 879 -42 0 FreeSans 80 0 0 0 Sw7
flabel locali 733 -124 768 -92 0 FreeSans 80 0 0 0 Sw7
flabel space 623 -126 658 -94 0 FreeSans 80 0 0 0 Sw6
flabel space 565 -124 600 -92 0 FreeSans 80 0 0 0 Sw5
flabel locali 456 -26 491 6 0 FreeSans 80 0 0 0 Sw4
flabel space 353 -10 388 22 0 FreeSans 80 0 0 0 Sw3
flabel space 289 -9 324 23 0 FreeSans 80 0 0 0 Sw2
flabel locali 204 -13 239 22 0 FreeSans 80 0 0 0 Sw1
flabel space 105 -25 147 17 0 FreeSans 80 0 0 0 Sw0
flabel locali -65 166 -41 187 0 FreeSans 80 0 0 0 vref_h
flabel metal1 -251 266 -207 304 0 FreeSans 80 0 0 0 vref_l
flabel locali -472 472 -421 523 0 FreeSans 80 0 0 0 samp_en
flabel space 6355 1428 6429 1499 0 FreeSans 80 0 0 0 Vout
<< properties >>
string FIXED_BBOX -193 -120 47 120
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 2.00 l 2.00 val 9.52 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

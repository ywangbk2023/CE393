** sch_path: /home/lcg3895/CE393/opamp_lna/low_noise_amp_tb_4.sch
**.subckt low_noise_amp_tb_4
x1 VDD net1 Vin_P Vin_N V0_P V0_N GND net1 Vbias Vref low_noise_amp
Vdd VDD GND 1.8
V2 Vbias GND 0.69
V3 Vref GND 0.35
VSource Vin_P Vin_N ac 1 sin(0 0.001 3000)
XC1 Vin_N V0_N sky130_fd_pr__cap_mim_m3_2 W=50 L=30 MF=1 m=1
XC2 Vin_P V0_P sky130_fd_pr__cap_mim_m3_2 W=50 L=30 MF=1 m=1
x3 VDD net2 V0_P V0_N V1_P V1_N GND net2 Vbias Vref low_noise_amp
x7 VDD net3 V1_P V1_N Vout_P Vout_N GND net3 Vbias Vref low_noise_amp
XC7 V1_N Vout_N sky130_fd_pr__cap_mim_m3_2 W=120 L=50 MF=1 m=1
XC6 V1_P Vout_P sky130_fd_pr__cap_mim_m3_2 W=120 L=50 MF=1 m=1
XC4 V0_N V1_N sky130_fd_pr__cap_mim_m3_2 W=75 L=30 MF=1 m=1
XC5 V0_P V1_P sky130_fd_pr__cap_mim_m3_2 W=75 L=30 MF=1 m=1
x2 Vin_P V0_P pseudoresistor
x4 Vin_N V0_N pseudoresistor
x5 V0_N V1_N pseudoresistor
x6 V0_P V1_P pseudoresistor
x8 V1_P Vout_P pseudoresistor
x9 V1_N Vout_N pseudoresistor
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ece393/open_pdks/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/ece393/open_pdks/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice



.PARAM R=0
.include postlayout_lna_extract.spice
.control
#noise v(Vout_P) Vsource dec 10 0.5 2000
tran 5us 1s
plot Vin_P-Vin_N Vout_P-Vout_N
#ac dec 10 0.000001 10000000
#plot vdb(V0_P) vdb(V0_N)
#plot vdb(V1_P) vdb(V1_N)
#plot vdb(Vout_P) vdb(Vout_N)
#plot vdb(V0_P) vdb(Vout_P)
save all
.endc

**** end user architecture code
**.ends

* expanding   symbol:  low_noise_amp.sym # of pins=10
** sym_path: /home/lcg3895/CE393/opamp_lna/low_noise_amp.sym
** sch_path: /home/lcg3895/CE393/opamp_lna/low_noise_amp.sch
.subckt low_noise_amp VDD Vcm_in INN INP V1P V1N VSS Vcm_out Vbias Vref
*.iopin VDD
*.iopin VSS
*.iopin Vbias
*.ipin INP
*.ipin INN
*.iopin Vref
*.iopin Vcm_in
*.iopin Vcm_out
*.opin V1N
*.opin V1P
XM3 CMFB Vref A0 VDD sky130_fd_pr__pfet_01v8 L=0.8 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 A0 Vbias VDD VDD sky130_fd_pr__pfet_01v8 L=0.8 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 V1N INP B0 VDD sky130_fd_pr__pfet_01v8 L=2 W=18 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 V1P INN B0 VDD sky130_fd_pr__pfet_01v8 L=2 W=18 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 V1N INP B1 VSS sky130_fd_pr__nfet_01v8 L=1 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 B0 Vbias VDD VDD sky130_fd_pr__pfet_01v8 L=0.8 W=4 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM13 B1 CMFB VSS VSS sky130_fd_pr__nfet_01v8 L=0.8 W=2 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM15 Vcm_out Vcm_out net1 Vcm_out sky130_fd_pr__pfet_01v8 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM16 net1 V1P V1P V1P sky130_fd_pr__pfet_01v8 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XM17 Vcm_out Vcm_out net2 Vcm_out sky130_fd_pr__pfet_01v8 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=5 m=5
XM18 net2 V1N V1N V1N sky130_fd_pr__pfet_01v8 L=0.6 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
XC1 Vcm_out VSS sky130_fd_pr__cap_mim_m3_1 W=0.1 L=0.1 MF=1 m=1
XM1 V1P INN B1 VSS sky130_fd_pr__nfet_01v8 L=1 W=12 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 A1 A1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.8 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 CMFB A1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.8 W=6 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 A1 Vcm_in A0 VDD sky130_fd_pr__pfet_01v8 L=0.8 W=8 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  /home/lcg3895/CE393/pseudoresistor.sym # of pins=2
** sym_path: /home/lcg3895/CE393/pseudoresistor.sym
** sch_path: /home/lcg3895/CE393/pseudoresistor.sch
.subckt pseudoresistor IN OUT
*.iopin IN
*.iopin OUT
XM5 net1 IN IN IN sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net2 net2 net1 net2 sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net3 net2 net2 net2 sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 OUT OUT net3 OUT sky130_fd_pr__pfet_01v8 L=0.5 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end

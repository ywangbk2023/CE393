magic
tech sky130A
magscale 1 2
timestamp 1701403287
<< nwell >>
rect -109 -662 109 662
<< pmos >>
rect -15 -600 15 600
<< pdiff >>
rect -73 588 -15 600
rect -73 -588 -61 588
rect -27 -588 -15 588
rect -73 -600 -15 -588
rect 15 588 73 600
rect 15 -588 27 588
rect 61 -588 73 588
rect 15 -600 73 -588
<< pdiffc >>
rect -61 -588 -27 588
rect 27 -588 61 588
<< poly >>
rect -15 600 15 626
rect -15 -626 15 -600
<< locali >>
rect -61 588 -27 604
rect -61 -604 -27 -588
rect 27 588 61 604
rect 27 -604 61 -588
<< viali >>
rect -61 -588 -27 588
rect 27 -588 61 588
<< metal1 >>
rect -67 588 -21 600
rect -67 -588 -61 588
rect -27 -588 -21 588
rect -67 -600 -21 -588
rect 21 588 67 600
rect 21 -588 27 588
rect 61 -588 67 588
rect 21 -600 67 -588
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 6 l 0.15 m 1 nf 1 diffcov 100 polycov 50 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

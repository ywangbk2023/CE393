magic
tech sky130A
magscale 1 2
timestamp 1701478054
<< nwell >>
rect -129 -249 129 249
<< pmos >>
rect -35 -187 35 187
<< pdiff >>
rect -93 175 -35 187
rect -93 -175 -81 175
rect -47 -175 -35 175
rect -93 -187 -35 -175
rect 35 175 93 187
rect 35 -175 47 175
rect 81 -175 93 175
rect 35 -187 93 -175
<< pdiffc >>
rect -81 -175 -47 175
rect 47 -175 81 175
<< poly >>
rect -35 187 35 213
rect -35 -213 35 -187
<< locali >>
rect -81 175 -47 191
rect -81 -191 -47 -175
rect 47 175 81 191
rect 47 -191 81 -175
<< viali >>
rect -81 -175 -47 175
rect 47 -175 81 175
<< metal1 >>
rect -87 175 -41 187
rect -87 -175 -81 175
rect -47 -175 -41 175
rect -87 -187 -41 -175
rect 41 175 87 187
rect 41 -175 47 175
rect 81 -175 87 175
rect 41 -187 87 -175
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.865 l 0.35 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1702102630
<< error_p >>
rect -29 132 29 138
rect -29 98 -17 132
rect -29 92 29 98
rect -29 -98 29 -92
rect -29 -132 -17 -98
rect -29 -138 29 -132
<< pwell >>
rect -211 -270 211 270
<< nmos >>
rect -15 -60 15 60
<< ndiff >>
rect -73 48 -15 60
rect -73 -48 -61 48
rect -27 -48 -15 48
rect -73 -60 -15 -48
rect 15 48 73 60
rect 15 -48 27 48
rect 61 -48 73 48
rect 15 -60 73 -48
<< ndiffc >>
rect -61 -48 -27 48
rect 27 -48 61 48
<< psubdiff >>
rect -175 200 -79 234
rect 79 200 175 234
rect -175 138 -141 200
rect 141 138 175 200
rect -175 -200 -141 -138
rect 141 -200 175 -138
rect -175 -234 -79 -200
rect 79 -234 175 -200
<< psubdiffcont >>
rect -79 200 79 234
rect -175 -138 -141 138
rect 141 -138 175 138
rect -79 -234 79 -200
<< poly >>
rect -33 132 33 148
rect -33 98 -17 132
rect 17 98 33 132
rect -33 82 33 98
rect -15 60 15 82
rect -15 -82 15 -60
rect -33 -98 33 -82
rect -33 -132 -17 -98
rect 17 -132 33 -98
rect -33 -148 33 -132
<< polycont >>
rect -17 98 17 132
rect -17 -132 17 -98
<< locali >>
rect -175 200 -79 234
rect 79 200 175 234
rect -175 138 -141 200
rect 141 138 175 200
rect -33 98 -17 132
rect 17 98 33 132
rect -61 48 -27 64
rect -61 -64 -27 -48
rect 27 48 61 64
rect 27 -64 61 -48
rect -33 -132 -17 -98
rect 17 -132 33 -98
rect -175 -200 -141 -138
rect 141 -200 175 -138
rect -175 -234 -79 -200
rect 79 -234 175 -200
<< viali >>
rect -17 98 17 132
rect -61 -48 -27 48
rect 27 -48 61 48
rect -17 -132 17 -98
<< metal1 >>
rect -29 132 29 138
rect -29 98 -17 132
rect 17 98 29 132
rect -29 92 29 98
rect -67 48 -21 60
rect -67 -48 -61 48
rect -27 -48 -21 48
rect -67 -60 -21 -48
rect 21 48 67 60
rect 21 -48 27 48
rect 61 -48 67 48
rect 21 -60 67 -48
rect -29 -98 29 -92
rect -29 -132 -17 -98
rect 17 -132 29 -98
rect -29 -138 29 -132
<< properties >>
string FIXED_BBOX -158 -217 158 217
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.6 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
timestamp 1702085311
<< nwell >>
rect -77 -81 77 81
<< pmos >>
rect -30 -50 30 50
<< pdiff >>
rect -59 44 -30 50
rect -59 -44 -53 44
rect -36 -44 -30 44
rect -59 -50 -30 -44
rect 30 44 59 50
rect 30 -44 36 44
rect 53 -44 59 44
rect 30 -50 59 -44
<< pdiffc >>
rect -53 -44 -36 44
rect 36 -44 53 44
<< poly >>
rect -30 50 30 63
rect -30 -63 30 -50
<< locali >>
rect -53 44 -36 52
rect -53 -52 -36 -44
rect 36 44 53 52
rect 36 -52 53 -44
<< viali >>
rect -53 -44 -36 44
rect 36 -44 53 44
<< metal1 >>
rect -56 44 -33 50
rect -56 -44 -53 44
rect -36 -44 -33 44
rect -56 -50 -33 -44
rect 33 44 56 50
rect 33 -44 36 44
rect 53 -44 56 44
rect 33 -50 56 -44
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.6 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
timestamp 1701908128
<< nwell >>
rect -276 -81 276 81
<< pmos >>
rect -229 -50 -179 50
rect -93 -50 -43 50
rect 43 -50 93 50
rect 179 -50 229 50
<< pdiff >>
rect -258 44 -229 50
rect -258 -44 -252 44
rect -235 -44 -229 44
rect -258 -50 -229 -44
rect -179 44 -150 50
rect -179 -44 -173 44
rect -156 -44 -150 44
rect -179 -50 -150 -44
rect -122 44 -93 50
rect -122 -44 -116 44
rect -99 -44 -93 44
rect -122 -50 -93 -44
rect -43 44 -14 50
rect -43 -44 -37 44
rect -20 -44 -14 44
rect -43 -50 -14 -44
rect 14 44 43 50
rect 14 -44 20 44
rect 37 -44 43 44
rect 14 -50 43 -44
rect 93 44 122 50
rect 93 -44 99 44
rect 116 -44 122 44
rect 93 -50 122 -44
rect 150 44 179 50
rect 150 -44 156 44
rect 173 -44 179 44
rect 150 -50 179 -44
rect 229 44 258 50
rect 229 -44 235 44
rect 252 -44 258 44
rect 229 -50 258 -44
<< pdiffc >>
rect -252 -44 -235 44
rect -173 -44 -156 44
rect -116 -44 -99 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 99 -44 116 44
rect 156 -44 173 44
rect 235 -44 252 44
<< poly >>
rect -229 50 -179 63
rect -93 50 -43 63
rect 43 50 93 63
rect 179 50 229 63
rect -229 -63 -179 -50
rect -93 -63 -43 -50
rect 43 -63 93 -50
rect 179 -63 229 -50
<< locali >>
rect -252 44 -235 52
rect -252 -52 -235 -44
rect -173 44 -156 52
rect -173 -52 -156 -44
rect -116 44 -99 52
rect -116 -52 -99 -44
rect -37 44 -20 52
rect -37 -52 -20 -44
rect 20 44 37 52
rect 20 -52 37 -44
rect 99 44 116 52
rect 99 -52 116 -44
rect 156 44 173 52
rect 156 -52 173 -44
rect 235 44 252 52
rect 235 -52 252 -44
<< viali >>
rect -252 -44 -235 44
rect -173 -44 -156 44
rect -116 -44 -99 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 99 -44 116 44
rect 156 -44 173 44
rect 235 -44 252 44
<< metal1 >>
rect -255 44 -232 50
rect -255 -44 -252 44
rect -235 -44 -232 44
rect -255 -50 -232 -44
rect -176 44 -153 50
rect -176 -44 -173 44
rect -156 -44 -153 44
rect -176 -50 -153 -44
rect -119 44 -96 50
rect -119 -44 -116 44
rect -99 -44 -96 44
rect -119 -50 -96 -44
rect -40 44 -17 50
rect -40 -44 -37 44
rect -20 -44 -17 44
rect -40 -50 -17 -44
rect 17 44 40 50
rect 17 -44 20 44
rect 37 -44 40 44
rect 17 -50 40 -44
rect 96 44 119 50
rect 96 -44 99 44
rect 116 -44 119 44
rect 96 -50 119 -44
rect 153 44 176 50
rect 153 -44 156 44
rect 173 -44 176 44
rect 153 -50 176 -44
rect 232 44 255 50
rect 232 -44 235 44
rect 252 -44 255 44
rect 232 -50 255 -44
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

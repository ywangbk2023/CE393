magic
tech sky130A
magscale 1 2
timestamp 1702102630
<< nwell >>
rect -186 -330 -88 -228
rect 92 -370 360 -76
rect 446 -394 644 -372
rect 446 -402 556 -394
rect 1294 -410 1548 -370
rect 814 -530 1118 -518
rect 814 -552 884 -530
rect 1054 -552 1118 -530
<< psubdiff >>
rect 20 -1278 118 -1254
rect 20 -1402 118 -1378
<< psubdiffcont >>
rect 20 -1378 118 -1278
<< poly >>
rect 1566 -356 1654 -334
rect 1566 -370 1606 -356
rect 446 -402 644 -372
rect 1294 -392 1606 -370
rect 1640 -392 1654 -356
rect 446 -490 562 -402
rect 1294 -410 1654 -392
rect 1566 -428 1654 -410
rect 444 -516 594 -490
rect 444 -602 466 -516
rect 548 -602 594 -516
rect 444 -652 594 -602
rect 814 -580 884 -528
rect 1054 -550 1124 -512
rect 1050 -580 1294 -550
rect 814 -688 858 -580
rect 642 -700 858 -688
rect 642 -708 808 -700
rect 550 -718 808 -708
rect 550 -738 674 -718
rect 550 -772 582 -738
rect 464 -788 582 -772
rect 642 -788 674 -738
rect 790 -734 808 -718
rect 842 -716 858 -700
rect 902 -638 992 -622
rect 902 -672 926 -638
rect 960 -672 992 -638
rect 902 -682 992 -672
rect 842 -734 860 -716
rect 790 -748 860 -734
rect 464 -803 674 -788
rect 224 -890 288 -874
rect 224 -924 238 -890
rect 272 -892 288 -890
rect 272 -922 408 -892
rect 272 -924 288 -922
rect 224 -942 288 -924
rect 464 -944 494 -803
rect 550 -816 674 -803
rect 902 -1112 932 -682
rect 1262 -796 1294 -580
rect 1010 -832 1294 -796
rect 1460 -790 1536 -774
rect 1460 -806 1480 -790
rect 1350 -830 1480 -806
rect 1524 -830 1536 -790
rect 1010 -846 1122 -832
rect 1350 -836 1536 -830
rect 1460 -846 1536 -836
rect 1010 -908 1036 -846
rect 1098 -908 1122 -846
rect 1010 -938 1122 -908
<< polycont >>
rect 1606 -392 1640 -356
rect 466 -602 548 -516
rect 582 -788 642 -738
rect 808 -734 842 -700
rect 926 -672 960 -638
rect 238 -924 272 -890
rect 1480 -830 1524 -790
rect 1036 -908 1098 -846
<< locali >>
rect 528 -134 562 -70
rect 896 -136 930 -66
rect 1008 -134 1042 -66
rect 1376 -134 1410 -70
rect 1168 -358 1250 -318
rect 1576 -354 1664 -334
rect 400 -374 434 -358
rect 338 -408 434 -374
rect 338 -808 372 -408
rect 414 -516 604 -458
rect 414 -602 466 -516
rect 548 -602 604 -516
rect 656 -514 690 -358
rect 1504 -426 1538 -356
rect 1304 -460 1538 -426
rect 1576 -406 1596 -354
rect 1642 -406 1664 -354
rect 1576 -440 1664 -406
rect 656 -544 802 -514
rect 656 -570 804 -544
rect 414 -654 604 -602
rect 704 -582 804 -570
rect 704 -664 754 -582
rect 548 -738 680 -704
rect 548 -788 582 -738
rect 642 -788 680 -738
rect 338 -842 454 -808
rect 548 -820 680 -788
rect 218 -890 292 -874
rect 218 -924 238 -890
rect 272 -924 292 -890
rect 218 -942 292 -924
rect 418 -942 454 -842
rect 716 -866 754 -664
rect 908 -636 994 -616
rect 908 -638 928 -636
rect 908 -672 926 -638
rect 962 -670 994 -636
rect 960 -672 994 -670
rect 908 -682 994 -672
rect 790 -700 858 -698
rect 790 -734 808 -700
rect 842 -716 858 -700
rect 1136 -716 1170 -514
rect 842 -718 1170 -716
rect 842 -734 1252 -718
rect 790 -752 1252 -734
rect 790 -754 1154 -752
rect 1008 -846 1122 -822
rect 1008 -866 1036 -846
rect 506 -900 1036 -866
rect 506 -902 754 -900
rect 506 -940 540 -902
rect 1008 -908 1036 -900
rect 1098 -908 1122 -846
rect 1214 -856 1252 -752
rect 1304 -856 1338 -460
rect 1460 -790 1536 -774
rect 1460 -830 1480 -790
rect 1524 -830 1536 -790
rect 1460 -846 1536 -830
rect 1008 -936 1122 -908
rect 668 -1050 978 -1042
rect 1392 -1050 1426 -978
rect 326 -1150 362 -1050
rect 668 -1078 1426 -1050
rect 668 -1150 704 -1078
rect 944 -1090 1426 -1078
rect 944 -1118 978 -1090
rect 326 -1188 704 -1150
rect 868 -1184 880 -1150
rect 20 -1278 118 -1262
rect 856 -1304 890 -1238
rect 20 -1394 118 -1378
<< viali >>
rect 528 -70 562 -36
rect 896 -66 930 -32
rect 1008 -66 1042 -32
rect 1376 -70 1410 -36
rect 1648 -210 1686 -174
rect -178 -366 -144 -332
rect -68 -412 -16 -372
rect 1596 -356 1642 -354
rect 1596 -392 1606 -356
rect 1606 -392 1640 -356
rect 1640 -392 1642 -356
rect 1596 -406 1642 -392
rect 1818 -384 1860 -342
rect 590 -786 632 -744
rect 928 -638 962 -636
rect 928 -670 960 -638
rect 960 -670 962 -638
rect 852 -1358 898 -1304
<< metal1 >>
rect 44 -32 1624 -2
rect 44 -36 896 -32
rect 44 -70 528 -36
rect 562 -66 896 -36
rect 930 -66 1008 -32
rect 1042 -36 1624 -32
rect 1042 -66 1376 -36
rect 562 -70 1376 -66
rect 1410 -70 1624 -36
rect 44 -76 1624 -70
rect 44 -90 380 -76
rect 1636 -160 1702 -148
rect 1624 -162 1702 -160
rect 1624 -222 1636 -162
rect 1698 -222 1702 -162
rect 1624 -236 1702 -222
rect -204 -310 -124 -304
rect -204 -380 -198 -310
rect -126 -380 -124 -310
rect 1624 -334 1678 -236
rect 1574 -346 1678 -334
rect 1792 -320 1910 -312
rect -204 -390 -124 -380
rect -94 -354 12 -346
rect -94 -434 -82 -354
rect -2 -362 12 -354
rect 1574 -354 1652 -346
rect -2 -402 262 -362
rect -2 -434 12 -402
rect -94 -444 12 -434
rect -102 -1252 -8 -646
rect 222 -726 262 -402
rect 1574 -406 1596 -354
rect 1642 -406 1652 -354
rect 1574 -410 1652 -406
rect 1570 -428 1652 -410
rect 1792 -398 1804 -320
rect 1896 -398 1910 -320
rect 1792 -416 1910 -398
rect 1570 -450 1602 -428
rect 1560 -466 1602 -450
rect 1534 -478 1602 -466
rect 1534 -494 1588 -478
rect 446 -614 578 -502
rect 1534 -614 1568 -494
rect 446 -616 1568 -614
rect 494 -636 1568 -616
rect 494 -642 928 -636
rect 918 -670 928 -642
rect 962 -642 1568 -636
rect 962 -670 990 -642
rect 1046 -644 1568 -642
rect 918 -682 990 -670
rect 554 -726 672 -706
rect 220 -744 672 -726
rect 220 -766 590 -744
rect 554 -786 590 -766
rect 632 -786 672 -744
rect 554 -812 672 -786
rect 1692 -1226 1770 -612
rect -102 -1258 164 -1252
rect -134 -1282 164 -1258
rect -136 -1284 196 -1282
rect 1692 -1284 1772 -1226
rect -136 -1304 1772 -1284
rect -136 -1358 852 -1304
rect 898 -1358 1772 -1304
rect -136 -1370 1772 -1358
rect -136 -1372 196 -1370
rect -134 -1396 164 -1372
rect -8 -1408 164 -1396
<< via1 >>
rect 1636 -174 1698 -162
rect 1636 -210 1648 -174
rect 1648 -210 1686 -174
rect 1686 -210 1698 -174
rect 1636 -222 1698 -210
rect -198 -332 -126 -310
rect -198 -366 -178 -332
rect -178 -366 -144 -332
rect -144 -366 -126 -332
rect -198 -380 -126 -366
rect -82 -372 -2 -354
rect -82 -412 -68 -372
rect -68 -412 -16 -372
rect -16 -412 -2 -372
rect -82 -434 -2 -412
rect 1804 -342 1896 -320
rect 1804 -384 1818 -342
rect 1818 -384 1860 -342
rect 1860 -384 1896 -342
rect 1804 -398 1896 -384
<< metal2 >>
rect 1636 -162 1702 -148
rect 1698 -222 1702 -162
rect 1636 -236 1702 -222
rect -202 -310 -124 -304
rect -202 -380 -198 -310
rect -126 -380 -124 -310
rect 1792 -320 1910 -314
rect -202 -392 -124 -380
rect -94 -354 14 -342
rect -94 -434 -82 -354
rect -2 -434 14 -354
rect 1792 -398 1804 -320
rect 1896 -398 1910 -320
rect 1792 -416 1910 -398
rect -94 -450 14 -434
use sky130_fd_pr__nfet_01v8_5TZ6LE  sky130_fd_pr__nfet_01v8_5TZ6LE_0
timestamp 1701820234
transform 1 0 479 0 1 -1004
box -73 -86 73 86
use sky130_fd_pr__nfet_01v8_5TZ6LE  sky130_fd_pr__nfet_01v8_5TZ6LE_1
timestamp 1701820234
transform 1 0 391 0 1 -1004
box -73 -86 73 86
use sky130_fd_pr__nfet_01v8_5TZ6LE  sky130_fd_pr__nfet_01v8_5TZ6LE_2
timestamp 1701820234
transform 1 0 1365 0 1 -918
box -73 -86 73 86
use sky130_fd_pr__nfet_01v8_5TZ6LE  sky130_fd_pr__nfet_01v8_5TZ6LE_3
timestamp 1701820234
transform 1 0 1277 0 1 -918
box -73 -86 73 86
use sky130_fd_pr__nfet_01v8_5TZ6LE  sky130_fd_pr__nfet_01v8_5TZ6LE_4
timestamp 1701820234
transform -1 0 917 0 -1 -1178
box -73 -86 73 86
use sky130_fd_pr__pfet_01v8_XCJR5L  sky130_fd_pr__pfet_01v8_XCJR5L_0
timestamp 1701819382
transform 1 0 609 0 1 -246
box -129 -170 129 170
use sky130_fd_pr__pfet_01v8_XCJR5L  sky130_fd_pr__pfet_01v8_XCJR5L_1
timestamp 1701819382
transform 1 0 481 0 1 -246
box -129 -170 129 170
use sky130_fd_pr__pfet_01v8_XCJR5L  sky130_fd_pr__pfet_01v8_XCJR5L_2
timestamp 1701819382
transform 1 0 1329 0 1 -246
box -129 -170 129 170
use sky130_fd_pr__pfet_01v8_XCJR5L  sky130_fd_pr__pfet_01v8_XCJR5L_3
timestamp 1701819382
transform 1 0 1457 0 1 -246
box -129 -170 129 170
use sky130_fd_pr__pfet_01v8_XCZ6WP  sky130_fd_pr__pfet_01v8_XCZ6WP_0
timestamp 1701819382
transform 1 0 849 0 1 -325
box -129 -249 129 249
use sky130_fd_pr__pfet_01v8_XCZ6WP  sky130_fd_pr__pfet_01v8_XCZ6WP_1
timestamp 1701819382
transform 1 0 1089 0 1 -325
box -129 -249 129 249
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0 ece393/open_pdks/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697562905
transform -1 0 1898 0 1 -594
box -38 -48 314 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_1 ece393/open_pdks/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697562905
transform -1 0 60 0 1 -630
box -38 -48 314 592
<< labels >>
flabel metal2 1804 -398 1896 -320 0 FreeSans 320 0 0 0 Clk
port 0 nsew
flabel polycont 256 -908 256 -908 0 FreeSans 320 0 0 0 Vref
port 1 nsew
flabel polycont 1502 -810 1502 -810 0 FreeSans 320 0 0 0 Vmac
port 2 nsew
flabel metal1 692 -38 692 -38 0 FreeSans 320 0 0 0 VDD
port 5 nsew
flabel metal1 614 -1336 614 -1336 0 FreeSans 320 0 0 0 VSS
port 4 nsew
flabel via1 -164 -350 -164 -350 0 FreeSans 320 0 0 0 Updown
port 3 nsew
<< end >>

magic
tech sky130A
timestamp 1702104985
<< nwell >>
rect -230 -81 230 81
<< pmos >>
rect -183 -50 -133 50
rect -104 -50 -54 50
rect -25 -50 25 50
rect 54 -50 104 50
rect 133 -50 183 50
<< pdiff >>
rect -212 44 -183 50
rect -212 -44 -206 44
rect -189 -44 -183 44
rect -212 -50 -183 -44
rect -133 44 -104 50
rect -133 -44 -127 44
rect -110 -44 -104 44
rect -133 -50 -104 -44
rect -54 44 -25 50
rect -54 -44 -48 44
rect -31 -44 -25 44
rect -54 -50 -25 -44
rect 25 44 54 50
rect 25 -44 31 44
rect 48 -44 54 44
rect 25 -50 54 -44
rect 104 44 133 50
rect 104 -44 110 44
rect 127 -44 133 44
rect 104 -50 133 -44
rect 183 44 212 50
rect 183 -44 189 44
rect 206 -44 212 44
rect 183 -50 212 -44
<< pdiffc >>
rect -206 -44 -189 44
rect -127 -44 -110 44
rect -48 -44 -31 44
rect 31 -44 48 44
rect 110 -44 127 44
rect 189 -44 206 44
<< poly >>
rect -183 50 -133 63
rect -104 50 -54 63
rect -25 50 25 63
rect 54 50 104 63
rect 133 50 183 63
rect -183 -63 -133 -50
rect -104 -63 -54 -50
rect -25 -63 25 -50
rect 54 -63 104 -50
rect 133 -63 183 -50
<< locali >>
rect -206 44 -189 52
rect -206 -52 -189 -44
rect -127 44 -110 52
rect -127 -52 -110 -44
rect -48 44 -31 52
rect -48 -52 -31 -44
rect 31 44 48 52
rect 31 -52 48 -44
rect 110 44 127 52
rect 110 -52 127 -44
rect 189 44 206 52
rect 189 -52 206 -44
<< viali >>
rect -206 -44 -189 44
rect -127 -44 -110 44
rect -48 -44 -31 44
rect 31 -44 48 44
rect 110 -44 127 44
rect 189 -44 206 44
<< metal1 >>
rect -209 44 -186 50
rect -209 -44 -206 44
rect -189 -44 -186 44
rect -209 -50 -186 -44
rect -130 44 -107 50
rect -130 -44 -127 44
rect -110 -44 -107 44
rect -130 -50 -107 -44
rect -51 44 -28 50
rect -51 -44 -48 44
rect -31 -44 -28 44
rect -51 -50 -28 -44
rect 28 44 51 50
rect 28 -44 31 44
rect 48 -44 51 44
rect 28 -50 51 -44
rect 107 44 130 50
rect 107 -44 110 44
rect 127 -44 130 44
rect 107 -50 130 -44
rect 186 44 209 50
rect 186 -44 189 44
rect 206 -44 209 44
rect 186 -50 209 -44
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.5 m 1 nf 5 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1701908128
<< metal3 >>
rect -5492 3012 -120 3040
rect -5492 -3012 -204 3012
rect -140 -3012 -120 3012
rect -5492 -3040 -120 -3012
rect 120 3012 5492 3040
rect 120 -3012 5408 3012
rect 5472 -3012 5492 3012
rect 120 -3040 5492 -3012
<< via3 >>
rect -204 -3012 -140 3012
rect 5408 -3012 5472 3012
<< mimcap >>
rect -5452 2960 -452 3000
rect -5452 -2960 -5412 2960
rect -492 -2960 -452 2960
rect -5452 -3000 -452 -2960
rect 160 2960 5160 3000
rect 160 -2960 200 2960
rect 5120 -2960 5160 2960
rect 160 -3000 5160 -2960
<< mimcapcontact >>
rect -5412 -2960 -492 2960
rect 200 -2960 5120 2960
<< metal4 >>
rect -220 3012 -124 3028
rect -5413 2960 -491 2961
rect -5413 -2960 -5412 2960
rect -492 -2960 -491 2960
rect -5413 -2961 -491 -2960
rect -220 -3012 -204 3012
rect -140 -3012 -124 3012
rect 5392 3012 5488 3028
rect 199 2960 5121 2961
rect 199 -2960 200 2960
rect 5120 -2960 5121 2960
rect 199 -2961 5121 -2960
rect -220 -3028 -124 -3012
rect 5392 -3012 5408 3012
rect 5472 -3012 5488 3012
rect 5392 -3028 5488 -3012
<< properties >>
string FIXED_BBOX 120 -3040 5200 3040
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 25 l 30 val 1.52k carea 2.00 cperi 0.19 nx 2 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

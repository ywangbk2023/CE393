magic
tech sky130A
magscale 1 2
timestamp 1701310363
<< nwell >>
rect -396 -1819 396 1819
<< pmos >>
rect -200 -1600 200 1600
<< pdiff >>
rect -258 1588 -200 1600
rect -258 -1588 -246 1588
rect -212 -1588 -200 1588
rect -258 -1600 -200 -1588
rect 200 1588 258 1600
rect 200 -1588 212 1588
rect 246 -1588 258 1588
rect 200 -1600 258 -1588
<< pdiffc >>
rect -246 -1588 -212 1588
rect 212 -1588 246 1588
<< nsubdiff >>
rect -360 1749 -264 1783
rect 264 1749 360 1783
rect -360 1687 -326 1749
rect 326 1687 360 1749
rect -360 -1749 -326 -1687
rect 326 -1749 360 -1687
rect -360 -1783 -264 -1749
rect 264 -1783 360 -1749
<< nsubdiffcont >>
rect -264 1749 264 1783
rect -360 -1687 -326 1687
rect 326 -1687 360 1687
rect -264 -1783 264 -1749
<< poly >>
rect -200 1681 200 1697
rect -200 1647 -184 1681
rect 184 1647 200 1681
rect -200 1600 200 1647
rect -200 -1647 200 -1600
rect -200 -1681 -184 -1647
rect 184 -1681 200 -1647
rect -200 -1697 200 -1681
<< polycont >>
rect -184 1647 184 1681
rect -184 -1681 184 -1647
<< locali >>
rect -360 1749 -264 1783
rect 264 1749 360 1783
rect -360 1687 -326 1749
rect 326 1687 360 1749
rect -200 1647 -184 1681
rect 184 1647 200 1681
rect -246 1588 -212 1604
rect -246 -1604 -212 -1588
rect 212 1588 246 1604
rect 212 -1604 246 -1588
rect -200 -1681 -184 -1647
rect 184 -1681 200 -1647
rect -360 -1749 -326 -1687
rect 326 -1749 360 -1687
rect -360 -1783 -264 -1749
rect 264 -1783 360 -1749
<< viali >>
rect -184 1647 184 1681
rect -246 -1588 -212 1588
rect 212 -1588 246 1588
rect -184 -1681 184 -1647
<< metal1 >>
rect -196 1681 196 1687
rect -196 1647 -184 1681
rect 184 1647 196 1681
rect -196 1641 196 1647
rect -252 1588 -206 1600
rect -252 -1588 -246 1588
rect -212 -1588 -206 1588
rect -252 -1600 -206 -1588
rect 206 1588 252 1600
rect 206 -1588 212 1588
rect 246 -1588 252 1588
rect 206 -1600 252 -1588
rect -196 -1647 196 -1641
rect -196 -1681 -184 -1647
rect 184 -1681 196 -1647
rect -196 -1687 196 -1681
<< properties >>
string FIXED_BBOX -343 -1766 343 1766
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 16 l 2 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

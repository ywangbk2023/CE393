** sch_path: /home/krr2464/CE393project/8bitADC_SARLOGIC_pinout.sch
**.subckt 8bitADC_SARLOGIC_pinout cmp start rstb clk dout0 doutb0 VSS VDD dout1 dout2 dout3 dout4
*+ dout5 dout6 dout7 doutb1 doutb2 doutb3 doutb4 doutb5 doutb6 doutb7
*.ipin cmp
*.ipin start
*.ipin rstb
*.ipin clk
*.iopin dout0
*.iopin doutb0
*.iopin VSS
*.iopin VDD
*.iopin dout1
*.iopin dout2
*.iopin dout3
*.iopin dout4
*.iopin dout5
*.iopin dout6
*.iopin dout7
*.iopin doutb1
*.iopin doutb2
*.iopin doutb3
*.iopin doutb4
*.iopin doutb5
*.iopin doutb6
*.iopin doutb7
x18 cmp VSS VNB VPB VDD cmp1 sky130_fd_sc_hd__buf_1
x19 clk VSS VNB VPB VDD net17 sky130_fd_sc_hd__buf_1
x20 net1 VSS VNB VPB VDD net2 sky130_fd_sc_hd__buf_1
x21 rstb VSS VNB VPB VDD net1 sky130_fd_sc_hd__buf_1
x22 start VSS VNB VPB VDD net8 sky130_fd_sc_hd__buf_1
x2 clk_t net8 net2 VSS VNB VPB VDD q q1 sky130_fd_sc_hd__dfrbp_1
x9 clk_t q net2 VSS VNB VPB VDD net9 q2 sky130_fd_sc_hd__dfrbp_1
x10 clk_t net9 net2 VSS VNB VPB VDD net10 q3 sky130_fd_sc_hd__dfrbp_1
x11 clk_t net10 net2 VSS VNB VPB VDD net11 net4 sky130_fd_sc_hd__dfrbp_1
x12 clk_t net11 net2 VSS VNB VPB VDD net12 net3 sky130_fd_sc_hd__dfrbp_1
x14 clk_t net12 net2 VSS VNB VPB VDD net13 net5 sky130_fd_sc_hd__dfrbp_1
x15 clk_t net13 net2 VSS VNB VPB VDD net14 net6 sky130_fd_sc_hd__dfrbp_1
x16 clk_t net14 net2 VSS VNB VPB VDD net15 net7 sky130_fd_sc_hd__dfrbp_1
x17 clk_t net15 net2 VSS VNB VPB VDD net16 net18 sky130_fd_sc_hd__dfrbp_1
x23 net17 VSS VNB VPB VDD clk_t sky130_fd_sc_hd__inv_1
x13 dout6 cmp1 net2 q1 VSS VNB VPB VDD dout7 doutb7 sky130_fd_sc_hd__dfbbp_1
x1 dout5 cmp1 net2 q2 VSS VNB VPB VDD dout6 doutb6 sky130_fd_sc_hd__dfbbp_1
x3 dout4 cmp1 net2 q3 VSS VNB VPB VDD dout5 doutb5 sky130_fd_sc_hd__dfbbp_1
x4 dout3 cmp1 net2 net4 VSS VNB VPB VDD dout4 doutb4 sky130_fd_sc_hd__dfbbp_1
x5 dout2 cmp1 net2 net3 VSS VNB VPB VDD dout3 doutb3 sky130_fd_sc_hd__dfbbp_1
x6 dout1 cmp1 net2 net5 VSS VNB VPB VDD dout2 doutb2 sky130_fd_sc_hd__dfbbp_1
x7 dout0 cmp1 net2 net6 VSS VNB VPB VDD dout1 doutb1 sky130_fd_sc_hd__dfbbp_1
x8 net16 cmp1 net2 net7 VSS VNB VPB VDD dout0 doutb0 sky130_fd_sc_hd__dfbbp_1
Vdd5 VDD GND 1.8
V1 CLK GND PULSE(0 1.8 0 0.1ns 0.1ns 2.5ns 5ns)
V3 VSS GND 0
Vdd7 trigger GND PWL(0 0.6 20ns 0.6 20.00001ns 1.2 25ns 1.2 25.00001ns 0.6 )
Vdd8 rstb GND PWL(0 1.2 5ns 1.2 5.00001ns 0.6 15ns 0.6 15.00001ns 1.2 )
Vdd1 samp_en GND PWL(0 0.6 5ns 0.6 5.00001ns 1.2 15ns 1.2 15.00001ns 0.6 )
V2 cmp GND PULSE(0 1.8 1.25ns 0.1ns 0.1ns 2.5ns 5ns)
**** begin user architecture code

** opencircuitdesign pdks install
.lib /home/ece393/open_pdks/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include /home/ece393/open_pdks/share/pdk/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice



.tran  0.01ns 100ns



**** end user architecture code
**.ends
.GLOBAL GND
.end

magic
tech sky130A
timestamp 1701309268
<< nwell >>
rect -87 -231 87 231
<< pmos >>
rect -40 -200 40 200
<< pdiff >>
rect -69 194 -40 200
rect -69 -194 -63 194
rect -46 -194 -40 194
rect -69 -200 -40 -194
rect 40 194 69 200
rect 40 -194 46 194
rect 63 -194 69 194
rect 40 -200 69 -194
<< pdiffc >>
rect -63 -194 -46 194
rect 46 -194 63 194
<< poly >>
rect -40 200 40 213
rect -40 -213 40 -200
<< locali >>
rect -63 194 -46 202
rect -63 -202 -46 -194
rect 46 194 63 202
rect 46 -202 63 -194
<< viali >>
rect -63 -194 -46 194
rect 46 -194 63 194
<< metal1 >>
rect -66 194 -43 200
rect -66 -194 -63 194
rect -46 -194 -43 194
rect -66 -200 -43 -194
rect 43 194 66 200
rect 43 -194 46 194
rect 63 -194 66 194
rect 43 -200 66 -194
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 4 l 0.8 m 1 nf 1 diffcov 100 polycov 100 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 100 rlcov 100 topc 0 botc 0 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>

magic
tech sky130A
magscale 1 2
timestamp 1702165270
<< nwell >>
rect 2038 626 2076 666
rect 2322 612 2358 648
rect 4430 620 4468 660
rect 6922 554 6960 590
rect 118 -56 288 -54
rect 762 -56 1034 -54
rect 118 -374 142 -56
rect 118 -376 374 -374
rect 742 -376 786 -56
rect 742 -378 1042 -376
rect 1318 -560 1354 -524
rect 7386 -618 7434 -372
rect 7386 -624 7556 -618
rect 302 -1358 336 -1324
rect 2692 -1366 2726 -1330
rect 7480 -1356 7516 -1322
rect 7484 -1446 7506 -1418
<< pwell >>
rect 4974 -736 5020 -702
rect 7764 -764 7818 -704
<< locali >>
rect -224 -58 -130 -10
rect -224 -60 -184 -58
rect 430 -64 470 8
rect 9184 -52 9190 -14
rect 9230 -52 9242 -14
rect 9184 -62 9242 -52
rect 7746 -116 7754 -82
<< viali >>
rect 2038 626 2076 666
rect 2322 612 2358 648
rect 4430 620 4468 660
rect 4712 626 4746 662
rect 7108 606 7144 640
rect 9492 630 9528 666
rect -76 564 -42 598
rect 6922 554 6960 590
rect 9214 548 9250 586
rect -248 426 -212 462
rect 20 428 56 462
rect 348 434 384 468
rect 1874 428 1912 466
rect 2412 436 2448 472
rect 2740 434 2776 468
rect 4268 426 4306 460
rect 4800 430 4840 466
rect 5142 440 5178 476
rect 6660 428 6696 464
rect 7198 414 7232 448
rect 7530 438 7564 474
rect 9048 430 9084 468
rect -76 296 -36 332
rect -38 44 2 82
rect 664 62 702 100
rect 1030 74 1066 110
rect 3128 60 3166 100
rect 5246 62 5282 98
rect 7358 64 7396 100
rect 9470 52 9510 96
rect -434 -48 -396 -6
rect 208 -54 246 -18
rect 1404 2 1442 42
rect 856 -44 894 -8
rect 2842 -46 2878 -10
rect 4954 -48 4988 -14
rect 7080 -46 7114 -10
rect 9190 -52 9230 -10
rect 1118 -106 1154 -70
rect 3246 -100 3282 -66
rect 3512 -116 3548 -82
rect 5352 -96 5392 -58
rect 5630 -116 5664 -82
rect 7474 -98 7510 -60
rect 7754 -118 7790 -82
rect 662 -202 706 -164
rect 3542 -504 3586 -466
rect 5664 -496 5702 -460
rect 7484 -504 7522 -464
rect 1318 -560 1354 -524
rect 9218 -594 9252 -558
rect 3136 -666 3174 -628
rect 5266 -662 5304 -624
rect 7374 -668 7408 -632
rect 9492 -666 9534 -626
rect -692 -728 -654 -690
rect 740 -744 782 -706
rect 1132 -774 1168 -738
rect 2846 -750 2894 -710
rect 4974 -736 5020 -702
rect 3252 -774 3288 -738
rect 5364 -770 5402 -734
rect 7092 -744 7136 -708
rect 7772 -752 7806 -718
rect 460 -1238 496 -1202
rect 1982 -1244 2018 -1210
rect 2312 -1240 2356 -1200
rect 2850 -1232 2886 -1198
rect 4370 -1256 4404 -1222
rect 4696 -1230 4738 -1188
rect 5238 -1234 5276 -1198
rect 6746 -1254 6784 -1216
rect 7634 -1244 7674 -1202
rect 9154 -1236 9188 -1202
rect 9488 -1238 9528 -1196
rect 7100 -1286 7134 -1252
rect 14 -1380 50 -1344
rect 302 -1358 336 -1324
rect 2692 -1366 2726 -1330
rect 5086 -1364 5122 -1330
rect 7480 -1356 7516 -1322
rect 2412 -1432 2446 -1398
rect 7192 -1426 7226 -1390
<< metal1 >>
rect -324 798 -172 800
rect -566 768 -172 798
rect -566 666 -536 768
rect -438 702 -172 768
rect -438 666 -418 702
rect -324 700 -172 702
rect -566 642 -418 666
rect 2026 666 2088 674
rect 2026 626 2038 666
rect 2076 626 2088 666
rect 4412 660 4486 672
rect -82 602 -28 610
rect 2026 608 2088 626
rect 2308 648 2370 658
rect 2308 612 2322 648
rect 2358 612 2370 648
rect 4412 620 4430 660
rect 4468 620 4486 660
rect 4412 612 4486 620
rect 4686 666 4768 674
rect 4686 614 4700 666
rect 4756 614 4768 666
rect 2308 602 2370 612
rect 4686 606 4768 614
rect 4808 670 4846 674
rect 4808 632 7034 670
rect 7204 666 9552 674
rect -82 534 -28 550
rect 6 480 76 528
rect 340 496 420 526
rect -266 462 -190 480
rect -266 426 -248 462
rect -212 426 -190 462
rect -266 402 -190 426
rect 4 468 84 480
rect 4 416 16 468
rect 72 416 84 468
rect 340 428 344 496
rect 414 428 420 496
rect 1844 478 1934 494
rect 340 422 420 428
rect 1484 438 1572 460
rect 4 400 84 416
rect 6 398 76 400
rect 1484 386 1502 438
rect 1554 386 1572 438
rect 1844 414 1860 478
rect 1926 414 1934 478
rect 2382 484 2478 504
rect 2382 428 2396 484
rect 2462 428 2478 484
rect 2382 416 2478 428
rect 2730 498 2810 530
rect 4808 510 4846 632
rect 6900 590 6968 602
rect 6900 554 6922 590
rect 6960 554 6968 590
rect 6900 542 6968 554
rect 2730 428 2732 498
rect 4238 490 4332 496
rect 2730 422 2810 428
rect 3870 426 3964 444
rect 1844 402 1934 414
rect 1484 364 1572 386
rect 3870 374 3886 426
rect 3940 374 3964 426
rect 4238 420 4250 490
rect 4326 420 4332 490
rect 4238 412 4332 420
rect 4790 466 4866 510
rect 4790 430 4800 466
rect 4840 430 4866 466
rect 4790 404 4866 430
rect 5122 500 5204 532
rect 7006 524 7034 632
rect 7082 664 7170 666
rect 7082 612 7088 664
rect 7158 612 7170 664
rect 7204 638 9492 666
rect 7082 606 7108 612
rect 7144 606 7170 612
rect 7082 568 7170 606
rect 7206 524 7240 638
rect 9486 630 9492 638
rect 9528 630 9552 666
rect 9486 612 9552 630
rect 9198 586 9274 598
rect 9198 548 9214 586
rect 9250 548 9274 586
rect 9198 534 9274 548
rect 5122 434 5128 500
rect 5198 434 5204 500
rect 6624 496 6726 510
rect 5122 424 5204 434
rect 6262 428 6358 448
rect 3870 360 3964 374
rect 6262 372 6278 428
rect 6342 372 6358 428
rect 6624 428 6636 496
rect 6714 428 6726 496
rect 7006 490 7244 524
rect 7514 500 7596 530
rect 6624 418 6726 428
rect 7180 460 7250 462
rect 7180 408 7190 460
rect 7244 408 7250 460
rect 7514 436 7522 500
rect 7588 436 7596 500
rect 9016 488 9112 494
rect 7514 424 7596 436
rect 8654 424 8738 442
rect 7180 398 7250 408
rect 6262 364 6358 372
rect 8654 370 8668 424
rect 8724 370 8738 424
rect 9016 414 9026 488
rect 9098 414 9112 488
rect 9016 408 9112 414
rect 8654 362 8738 370
rect -88 354 -14 360
rect -88 290 -82 354
rect -16 290 -14 354
rect -88 282 -14 290
rect -568 158 -334 254
rect 26 160 784 256
rect -568 -162 -472 158
rect 652 126 730 128
rect -64 92 14 124
rect -64 36 -56 92
rect 8 36 14 92
rect 650 118 736 126
rect 650 48 656 118
rect 730 48 736 118
rect 1020 110 1078 126
rect 1014 106 1030 110
rect 1066 106 1084 110
rect 1014 54 1022 106
rect 1074 54 1084 106
rect 3112 102 3198 124
rect 1014 48 1084 54
rect 1374 56 1468 94
rect 650 40 736 48
rect -64 28 14 36
rect -444 -6 -376 8
rect -444 -48 -434 -6
rect -396 -48 -376 -6
rect -444 -66 -376 -48
rect 196 -18 260 -2
rect 196 -54 208 -18
rect 246 -54 260 -18
rect 196 -64 260 -54
rect 834 -8 904 6
rect 834 -44 856 -8
rect 894 -44 904 -8
rect 1374 -10 1388 56
rect 1458 -10 1468 56
rect 1374 -20 1468 -10
rect 2480 46 2592 76
rect 3112 50 3128 102
rect 3186 50 3198 102
rect 5222 110 5314 126
rect 3112 46 3198 50
rect 2480 -32 2498 46
rect 2586 -32 2592 46
rect 4586 36 4704 62
rect 5222 52 5238 110
rect 5292 52 5314 110
rect 7338 112 7432 128
rect 7338 56 7352 112
rect 7416 56 7432 112
rect 9454 110 9536 122
rect 5222 44 5314 52
rect 1106 -42 1170 -40
rect 834 -62 904 -44
rect 1096 -52 1170 -42
rect 2480 -46 2592 -32
rect 2812 -10 2906 18
rect 2812 -46 2842 -10
rect 2878 -46 2906 -10
rect 4586 -44 4608 36
rect 4686 -44 4704 36
rect 6724 36 6814 52
rect 7338 42 7432 56
rect 1096 -114 1102 -52
rect 1164 -114 1170 -52
rect 2812 -66 2906 -46
rect 1096 -120 1170 -114
rect 1106 -122 1170 -120
rect -1166 -258 -472 -162
rect 648 -144 740 -138
rect 648 -222 662 -144
rect 736 -222 740 -144
rect 2826 -156 2882 -66
rect 3204 -114 3210 -46
rect 3278 -66 3290 -46
rect 4586 -58 4704 -44
rect 4938 -14 5012 12
rect 4938 -48 4954 -14
rect 4988 -48 5012 -14
rect 6724 -34 6738 36
rect 6804 -34 6814 36
rect 8840 38 8946 60
rect 4938 -60 5012 -48
rect 5306 -46 5398 -34
rect 3282 -100 3290 -66
rect 3490 -82 3572 -76
rect 3490 -84 3512 -82
rect 3278 -114 3290 -100
rect 3204 -120 3290 -114
rect 3336 -114 3512 -84
rect 3336 -156 3368 -114
rect 3490 -116 3512 -114
rect 3548 -116 3572 -82
rect 3490 -122 3572 -116
rect 2826 -190 3368 -156
rect 4962 -162 4990 -60
rect 5306 -116 5316 -46
rect 5394 -116 5398 -46
rect 6724 -52 6814 -34
rect 7066 -10 7126 0
rect 7066 -46 7080 -10
rect 7114 -46 7126 -10
rect 7066 -54 7126 -46
rect 7414 -36 7520 -24
rect 5612 -82 5678 -74
rect 5612 -84 5630 -82
rect 5306 -122 5398 -116
rect 5448 -112 5630 -84
rect 5448 -162 5478 -112
rect 5612 -116 5630 -112
rect 5664 -116 5678 -82
rect 5612 -126 5678 -116
rect 4962 -190 5478 -162
rect 7080 -172 7108 -54
rect 7414 -112 7430 -36
rect 7502 -60 7520 -36
rect 8840 -36 8860 38
rect 8932 -36 8946 38
rect 9454 46 9466 110
rect 9524 46 9536 110
rect 9454 36 9536 46
rect 8840 -50 8946 -36
rect 9172 -10 9244 6
rect 7510 -98 7520 -60
rect 9172 -52 9190 -10
rect 9230 -52 9244 -10
rect 7736 -82 7804 -74
rect 7736 -84 7754 -82
rect 7502 -112 7520 -98
rect 7414 -122 7520 -112
rect 7570 -114 7754 -84
rect 7570 -172 7598 -114
rect 7736 -118 7754 -114
rect 7790 -118 7804 -82
rect 7736 -124 7804 -118
rect 9172 -158 9244 -52
rect 7080 -200 7598 -172
rect 9170 -198 9646 -158
rect 648 -230 740 -222
rect -1165 -835 -1071 -258
rect -300 -308 -174 -278
rect -300 -372 -274 -308
rect -206 -372 -174 -308
rect -300 -400 -174 -372
rect 3502 -452 3618 -432
rect 1282 -504 1392 -494
rect 1282 -572 1302 -504
rect 1384 -572 1392 -504
rect 3502 -514 3516 -452
rect 3600 -514 3618 -452
rect 3502 -526 3618 -514
rect 5630 -444 5734 -424
rect 5630 -508 5646 -444
rect 5720 -508 5734 -444
rect 5630 -530 5734 -508
rect 7456 -454 7566 -424
rect 9608 -434 9646 -198
rect 7456 -514 7480 -454
rect 7548 -514 7566 -454
rect 9404 -470 9646 -434
rect 7456 -530 7566 -514
rect 1282 -586 1392 -572
rect 9178 -558 9280 -550
rect 1012 -620 1090 -606
rect -722 -680 -618 -662
rect 1012 -672 1024 -620
rect 1076 -672 1090 -620
rect 3128 -618 3214 -602
rect 1012 -680 1090 -672
rect 1724 -652 1812 -626
rect -722 -734 -702 -680
rect -630 -734 -618 -680
rect -722 -752 -618 -734
rect 222 -698 344 -686
rect 222 -760 238 -698
rect 338 -760 344 -698
rect 222 -770 344 -760
rect 710 -704 828 -692
rect 710 -780 726 -704
rect 810 -780 828 -704
rect 710 -800 828 -780
rect 1122 -726 1234 -708
rect 1122 -738 1138 -726
rect 1122 -774 1132 -738
rect 1122 -786 1138 -774
rect 1208 -786 1234 -726
rect 1724 -710 1746 -652
rect 1808 -710 1812 -652
rect 3128 -628 3146 -618
rect 3128 -666 3136 -628
rect 3128 -670 3146 -666
rect 3198 -670 3214 -618
rect 5246 -608 5326 -588
rect 3128 -684 3214 -670
rect 3844 -644 3934 -624
rect 1724 -728 1812 -710
rect 2832 -702 2948 -688
rect 2832 -764 2842 -702
rect 2928 -764 2948 -702
rect 2832 -780 2948 -764
rect 3240 -718 3356 -698
rect 3240 -738 3272 -718
rect 3240 -774 3252 -738
rect 3240 -780 3272 -774
rect 3336 -780 3356 -718
rect 3844 -716 3856 -644
rect 3924 -716 3934 -644
rect 5246 -662 5266 -608
rect 5320 -660 5326 -608
rect 7358 -608 7454 -584
rect 9178 -594 9218 -558
rect 9252 -560 9280 -558
rect 9402 -560 9442 -470
rect 9252 -562 9442 -560
rect 9252 -592 9440 -562
rect 9474 -578 9608 -552
rect 9252 -594 9280 -592
rect 9178 -602 9280 -594
rect 5304 -662 5326 -660
rect 5246 -676 5326 -662
rect 5960 -650 6044 -622
rect 3844 -726 3934 -716
rect 4930 -696 5060 -686
rect 1122 -802 1234 -786
rect 3240 -800 3356 -780
rect 4930 -762 4946 -696
rect 5046 -762 5060 -696
rect 4930 -784 5060 -762
rect 5356 -698 5486 -676
rect 5356 -734 5390 -698
rect 5356 -770 5364 -734
rect 5464 -768 5486 -698
rect 5960 -716 5970 -650
rect 6038 -716 6044 -650
rect 7358 -676 7372 -608
rect 7438 -676 7454 -608
rect 7358 -684 7454 -676
rect 8074 -644 8160 -628
rect 5960 -726 6044 -716
rect 7068 -708 7154 -696
rect 7068 -744 7092 -708
rect 7136 -722 7154 -708
rect 7764 -718 7818 -704
rect 7764 -722 7772 -718
rect 7136 -744 7772 -722
rect 7068 -752 7772 -744
rect 7806 -752 7818 -718
rect 8074 -714 8084 -644
rect 8152 -714 8160 -644
rect 9474 -678 9490 -578
rect 9586 -678 9608 -578
rect 9474 -690 9608 -678
rect 8074 -724 8160 -714
rect 7068 -758 7818 -752
rect 7068 -760 7154 -758
rect 7764 -764 7818 -758
rect 5402 -770 5486 -768
rect 5356 -790 5486 -770
rect -1165 -929 -915 -835
rect -294 -992 -186 -978
rect -294 -1072 -286 -992
rect -200 -1050 -186 -992
rect -200 -1072 -49 -1050
rect -294 -1080 -49 -1072
rect -79 -1231 -49 -1080
rect 8730 -1106 8832 -1090
rect 792 -1142 902 -1126
rect 434 -1184 528 -1174
rect -79 -1261 233 -1231
rect -14 -1332 82 -1310
rect -14 -1390 4 -1332
rect 66 -1390 82 -1332
rect -14 -1406 82 -1390
rect 6 -1428 66 -1406
rect 203 -1555 233 -1261
rect 434 -1254 442 -1184
rect 520 -1254 528 -1184
rect 792 -1200 810 -1142
rect 884 -1200 902 -1142
rect 1558 -1172 1638 -1108
rect 3228 -1136 3320 -1122
rect 2294 -1172 2400 -1150
rect 792 -1210 902 -1200
rect 1954 -1200 2030 -1194
rect 434 -1268 528 -1254
rect 1954 -1266 1962 -1200
rect 2028 -1266 2030 -1200
rect 1954 -1298 2030 -1266
rect 2294 -1246 2310 -1172
rect 2386 -1246 2400 -1172
rect 2294 -1268 2400 -1246
rect 2828 -1186 2920 -1184
rect 2828 -1246 2836 -1186
rect 2906 -1246 2920 -1186
rect 3228 -1194 3244 -1136
rect 3306 -1194 3320 -1136
rect 5576 -1142 5680 -1118
rect 4674 -1172 4774 -1154
rect 3228 -1206 3320 -1194
rect 2828 -1252 2920 -1246
rect 4344 -1214 4424 -1194
rect 4344 -1282 4356 -1214
rect 4422 -1282 4424 -1214
rect 4674 -1240 4690 -1172
rect 4760 -1240 4774 -1172
rect 4674 -1256 4774 -1240
rect 5218 -1182 5314 -1178
rect 5218 -1248 5226 -1182
rect 5294 -1248 5314 -1182
rect 5576 -1200 5594 -1142
rect 5664 -1200 5680 -1142
rect 7076 -1178 7198 -1150
rect 8730 -1162 8748 -1106
rect 8806 -1162 8832 -1106
rect 5576 -1210 5680 -1200
rect 6734 -1208 6816 -1196
rect 5218 -1254 5314 -1248
rect 4344 -1300 4424 -1282
rect 6734 -1276 6738 -1208
rect 6812 -1276 6816 -1208
rect 7076 -1252 7098 -1178
rect 7174 -1252 7198 -1178
rect 7076 -1274 7100 -1252
rect 6734 -1300 6816 -1276
rect 7080 -1286 7100 -1274
rect 7134 -1274 7198 -1252
rect 7616 -1184 7700 -1166
rect 8730 -1172 8832 -1162
rect 9498 -1170 9528 -1168
rect 7616 -1254 7622 -1184
rect 7694 -1254 7700 -1184
rect 7616 -1260 7700 -1254
rect 9130 -1202 9204 -1192
rect 9130 -1264 9136 -1202
rect 9198 -1264 9204 -1202
rect 7134 -1286 7150 -1274
rect 7080 -1298 7150 -1286
rect 9130 -1296 9204 -1264
rect 9474 -1196 9540 -1170
rect 9474 -1238 9488 -1196
rect 9528 -1238 9540 -1196
rect 9474 -1262 9540 -1238
rect 9474 -1296 9662 -1262
rect 288 -1324 354 -1314
rect 288 -1358 302 -1324
rect 336 -1358 354 -1324
rect 288 -1370 354 -1358
rect 2674 -1330 2746 -1312
rect 2674 -1366 2692 -1330
rect 2726 -1366 2746 -1330
rect 2674 -1376 2746 -1366
rect 4766 -1352 4876 -1324
rect 2392 -1384 2458 -1376
rect 2392 -1436 2398 -1384
rect 2452 -1436 2458 -1384
rect 4766 -1418 4784 -1352
rect 4854 -1418 4876 -1352
rect 5072 -1330 5140 -1316
rect 5072 -1364 5086 -1330
rect 5122 -1364 5140 -1330
rect 5072 -1376 5140 -1364
rect 7454 -1322 7540 -1296
rect 9474 -1302 9540 -1296
rect 7454 -1356 7480 -1322
rect 7516 -1356 7540 -1322
rect 7454 -1370 7540 -1356
rect 4766 -1436 4876 -1418
rect 7178 -1390 7244 -1380
rect 7178 -1426 7192 -1390
rect 7226 -1426 7244 -1390
rect 2392 -1442 2458 -1436
rect 7178 -1442 7244 -1426
rect 4678 -1606 7016 -1604
rect 4596 -1630 7016 -1606
rect 4596 -1636 6946 -1630
rect 4596 -1704 4628 -1636
rect 4708 -1644 6946 -1636
rect 4708 -1704 4736 -1644
rect 6938 -1682 6946 -1644
rect 7008 -1682 7016 -1630
rect 6938 -1686 7016 -1682
rect 7074 -1614 7176 -1612
rect 9624 -1614 9662 -1296
rect 7074 -1628 9662 -1614
rect 7074 -1682 7100 -1628
rect 7154 -1654 9662 -1628
rect 7154 -1682 7176 -1654
rect 7074 -1700 7176 -1682
rect 4596 -1740 4736 -1704
<< via1 >>
rect -536 666 -438 768
rect 4700 662 4756 666
rect 4700 626 4712 662
rect 4712 626 4746 662
rect 4746 626 4756 662
rect 4700 614 4756 626
rect -82 598 -28 602
rect -82 564 -76 598
rect -76 564 -42 598
rect -42 564 -28 598
rect -82 550 -28 564
rect 16 462 72 468
rect 16 428 20 462
rect 20 428 56 462
rect 56 428 72 462
rect 16 416 72 428
rect 344 468 414 496
rect 344 434 348 468
rect 348 434 384 468
rect 384 434 414 468
rect 344 428 414 434
rect 1502 386 1554 438
rect 1860 466 1926 478
rect 1860 428 1874 466
rect 1874 428 1912 466
rect 1912 428 1926 466
rect 1860 414 1926 428
rect 2396 472 2462 484
rect 2396 436 2412 472
rect 2412 436 2448 472
rect 2448 436 2462 472
rect 2396 428 2462 436
rect 2732 468 2810 498
rect 2732 434 2740 468
rect 2740 434 2776 468
rect 2776 434 2810 468
rect 2732 428 2810 434
rect 3886 374 3940 426
rect 4250 460 4326 490
rect 4250 426 4268 460
rect 4268 426 4306 460
rect 4306 426 4326 460
rect 4250 420 4326 426
rect 7088 640 7158 664
rect 7088 612 7108 640
rect 7108 612 7144 640
rect 7144 612 7158 640
rect 5128 476 5198 500
rect 5128 440 5142 476
rect 5142 440 5178 476
rect 5178 440 5198 476
rect 5128 434 5198 440
rect 6278 372 6342 428
rect 6636 464 6714 496
rect 6636 428 6660 464
rect 6660 428 6696 464
rect 6696 428 6714 464
rect 7190 448 7244 460
rect 7190 414 7198 448
rect 7198 414 7232 448
rect 7232 414 7244 448
rect 7190 408 7244 414
rect 7522 474 7588 500
rect 7522 438 7530 474
rect 7530 438 7564 474
rect 7564 438 7588 474
rect 7522 436 7588 438
rect 8668 370 8724 424
rect 9026 468 9098 488
rect 9026 430 9048 468
rect 9048 430 9084 468
rect 9084 430 9098 468
rect 9026 414 9098 430
rect -82 332 -16 354
rect -82 296 -76 332
rect -76 296 -36 332
rect -36 296 -16 332
rect -82 290 -16 296
rect -56 82 8 92
rect -56 44 -38 82
rect -38 44 2 82
rect 2 44 8 82
rect -56 36 8 44
rect 656 100 730 118
rect 656 62 664 100
rect 664 62 702 100
rect 702 62 730 100
rect 656 48 730 62
rect 1022 74 1030 106
rect 1030 74 1066 106
rect 1066 74 1074 106
rect 1022 54 1074 74
rect 1388 42 1458 56
rect 1388 2 1404 42
rect 1404 2 1442 42
rect 1442 2 1458 42
rect 1388 -10 1458 2
rect 3128 100 3186 102
rect 3128 60 3166 100
rect 3166 60 3186 100
rect 3128 50 3186 60
rect 2498 -32 2586 46
rect 5238 98 5292 110
rect 5238 62 5246 98
rect 5246 62 5282 98
rect 5282 62 5292 98
rect 5238 52 5292 62
rect 7352 100 7416 112
rect 7352 64 7358 100
rect 7358 64 7396 100
rect 7396 64 7416 100
rect 7352 56 7416 64
rect 4608 -44 4686 36
rect 1102 -70 1164 -52
rect 1102 -106 1118 -70
rect 1118 -106 1154 -70
rect 1154 -106 1164 -70
rect 1102 -114 1164 -106
rect 662 -164 736 -144
rect 662 -202 706 -164
rect 706 -202 736 -164
rect 662 -222 736 -202
rect 3210 -66 3278 -46
rect 6738 -34 6804 36
rect 3210 -100 3246 -66
rect 3246 -100 3278 -66
rect 3210 -114 3278 -100
rect 5316 -58 5394 -46
rect 5316 -96 5352 -58
rect 5352 -96 5392 -58
rect 5392 -96 5394 -58
rect 5316 -116 5394 -96
rect 7430 -60 7502 -36
rect 8860 -36 8932 38
rect 9466 96 9524 110
rect 9466 52 9470 96
rect 9470 52 9510 96
rect 9510 52 9524 96
rect 9466 46 9524 52
rect 7430 -98 7474 -60
rect 7474 -98 7502 -60
rect 7430 -112 7502 -98
rect -274 -372 -206 -308
rect 1302 -524 1384 -504
rect 1302 -560 1318 -524
rect 1318 -560 1354 -524
rect 1354 -560 1384 -524
rect 1302 -572 1384 -560
rect 3516 -466 3600 -452
rect 3516 -504 3542 -466
rect 3542 -504 3586 -466
rect 3586 -504 3600 -466
rect 3516 -514 3600 -504
rect 5646 -460 5720 -444
rect 5646 -496 5664 -460
rect 5664 -496 5702 -460
rect 5702 -496 5720 -460
rect 5646 -508 5720 -496
rect 7480 -464 7548 -454
rect 7480 -504 7484 -464
rect 7484 -504 7522 -464
rect 7522 -504 7548 -464
rect 7480 -514 7548 -504
rect 1024 -672 1076 -620
rect -702 -690 -630 -680
rect -702 -728 -692 -690
rect -692 -728 -654 -690
rect -654 -728 -630 -690
rect -702 -734 -630 -728
rect 238 -760 338 -698
rect 726 -706 810 -704
rect 726 -744 740 -706
rect 740 -744 782 -706
rect 782 -744 810 -706
rect 726 -780 810 -744
rect 1138 -738 1208 -726
rect 1138 -774 1168 -738
rect 1168 -774 1208 -738
rect 1138 -786 1208 -774
rect 1746 -710 1808 -652
rect 3146 -628 3198 -618
rect 3146 -666 3174 -628
rect 3174 -666 3198 -628
rect 3146 -670 3198 -666
rect 2842 -710 2928 -702
rect 2842 -750 2846 -710
rect 2846 -750 2894 -710
rect 2894 -750 2928 -710
rect 2842 -764 2928 -750
rect 3272 -738 3336 -718
rect 3272 -774 3288 -738
rect 3288 -774 3336 -738
rect 3272 -780 3336 -774
rect 3856 -716 3924 -644
rect 5266 -624 5320 -608
rect 5266 -660 5304 -624
rect 5304 -660 5320 -624
rect 4946 -702 5046 -696
rect 4946 -736 4974 -702
rect 4974 -736 5020 -702
rect 5020 -736 5046 -702
rect 4946 -762 5046 -736
rect 5390 -734 5464 -698
rect 5390 -768 5402 -734
rect 5402 -768 5464 -734
rect 5970 -716 6038 -650
rect 7372 -632 7438 -608
rect 7372 -668 7374 -632
rect 7374 -668 7408 -632
rect 7408 -668 7438 -632
rect 7372 -676 7438 -668
rect 8084 -714 8152 -644
rect 9490 -626 9586 -578
rect 9490 -666 9492 -626
rect 9492 -666 9534 -626
rect 9534 -666 9586 -626
rect 9490 -678 9586 -666
rect -286 -1072 -200 -992
rect 4 -1344 66 -1332
rect 4 -1380 14 -1344
rect 14 -1380 50 -1344
rect 50 -1380 66 -1344
rect 4 -1390 66 -1380
rect 442 -1202 520 -1184
rect 442 -1238 460 -1202
rect 460 -1238 496 -1202
rect 496 -1238 520 -1202
rect 442 -1254 520 -1238
rect 810 -1200 884 -1142
rect 1962 -1210 2028 -1200
rect 1962 -1244 1982 -1210
rect 1982 -1244 2018 -1210
rect 2018 -1244 2028 -1210
rect 1962 -1266 2028 -1244
rect 2310 -1200 2386 -1172
rect 2310 -1240 2312 -1200
rect 2312 -1240 2356 -1200
rect 2356 -1240 2386 -1200
rect 2310 -1246 2386 -1240
rect 2836 -1198 2906 -1186
rect 2836 -1232 2850 -1198
rect 2850 -1232 2886 -1198
rect 2886 -1232 2906 -1198
rect 2836 -1246 2906 -1232
rect 3244 -1194 3306 -1136
rect 4356 -1222 4422 -1214
rect 4356 -1256 4370 -1222
rect 4370 -1256 4404 -1222
rect 4404 -1256 4422 -1222
rect 4356 -1282 4422 -1256
rect 4690 -1188 4760 -1172
rect 4690 -1230 4696 -1188
rect 4696 -1230 4738 -1188
rect 4738 -1230 4760 -1188
rect 4690 -1240 4760 -1230
rect 5226 -1198 5294 -1182
rect 5226 -1234 5238 -1198
rect 5238 -1234 5276 -1198
rect 5276 -1234 5294 -1198
rect 5226 -1248 5294 -1234
rect 5594 -1200 5664 -1142
rect 8748 -1162 8806 -1106
rect 6738 -1216 6812 -1208
rect 6738 -1254 6746 -1216
rect 6746 -1254 6784 -1216
rect 6784 -1254 6812 -1216
rect 6738 -1276 6812 -1254
rect 7098 -1252 7174 -1178
rect 7622 -1202 7694 -1184
rect 7622 -1244 7634 -1202
rect 7634 -1244 7674 -1202
rect 7674 -1244 7694 -1202
rect 7622 -1254 7694 -1244
rect 9136 -1236 9154 -1202
rect 9154 -1236 9188 -1202
rect 9188 -1236 9198 -1202
rect 9136 -1264 9198 -1236
rect 2398 -1398 2452 -1384
rect 2398 -1432 2412 -1398
rect 2412 -1432 2446 -1398
rect 2446 -1432 2452 -1398
rect 2398 -1436 2452 -1432
rect 4784 -1418 4854 -1352
rect 4628 -1704 4708 -1636
rect 6946 -1682 7008 -1630
rect 7100 -1682 7154 -1628
<< metal2 >>
rect -566 768 -418 798
rect -566 666 -536 768
rect -438 666 -418 768
rect -566 642 -418 666
rect -146 726 4744 758
rect -146 448 -114 726
rect 4712 674 4744 726
rect 9544 705 9596 706
rect 7080 674 7174 686
rect 4688 666 4770 674
rect 4688 614 4700 666
rect 4756 614 4770 666
rect -82 602 -28 610
rect 4688 608 4770 614
rect 7080 612 7088 674
rect 7158 612 7174 674
rect 7080 606 7174 612
rect 8851 676 9596 705
rect 8851 675 9536 676
rect -28 550 7592 578
rect -82 534 -28 550
rect 340 496 420 550
rect 4 468 84 480
rect 4 448 16 468
rect -146 416 16 448
rect 72 416 84 468
rect 340 428 344 496
rect 414 428 420 496
rect 1844 478 1934 494
rect 340 422 420 428
rect 1484 448 1572 460
rect -16 414 84 416
rect 4 400 84 414
rect 1484 392 1500 448
rect 1558 392 1572 448
rect 1844 414 1860 478
rect 1926 414 1934 478
rect 2382 484 2478 504
rect 2382 428 2396 484
rect 2462 428 2478 484
rect 2382 416 2478 428
rect 2730 498 2810 550
rect 2730 428 2732 498
rect 5122 500 5204 550
rect 7514 530 7592 550
rect 4238 490 4332 496
rect 2730 422 2810 428
rect 3870 432 3964 444
rect 1844 402 1934 414
rect 1484 386 1502 392
rect 1554 386 1572 392
rect 1484 364 1572 386
rect -90 354 -10 362
rect -90 290 -82 354
rect -16 324 -10 354
rect 1872 332 1926 402
rect 3870 374 3886 432
rect 3944 374 3964 432
rect 4238 420 4250 490
rect 4326 420 4332 490
rect 5122 434 5128 500
rect 5198 434 5204 500
rect 6624 496 6726 510
rect 5122 424 5204 434
rect 6262 428 6358 448
rect 4238 412 4332 420
rect 3870 360 3964 374
rect 4268 332 4308 412
rect 6262 372 6278 428
rect 6342 372 6358 428
rect 6624 428 6636 496
rect 6714 428 6726 496
rect 7514 500 7596 530
rect 8851 505 8881 675
rect 6624 418 6726 428
rect 7180 460 7250 462
rect 6262 364 6358 372
rect 6660 332 6692 418
rect 7180 408 7190 460
rect 7244 428 7250 460
rect 7514 436 7522 500
rect 7588 436 7596 500
rect 7244 408 7483 428
rect 7514 424 7596 436
rect 8593 475 8881 505
rect 8935 543 9171 573
rect 7180 398 7483 408
rect 7453 391 7483 398
rect 8593 391 8623 475
rect 8935 442 8965 543
rect 7453 361 8623 391
rect 8654 424 8965 442
rect 8654 370 8668 424
rect 8724 412 8965 424
rect 9016 488 9112 494
rect 9016 414 9026 488
rect 9098 414 9112 488
rect 8724 370 8738 412
rect 9016 408 9112 414
rect 8654 362 8738 370
rect 9058 332 9100 408
rect -16 290 85 324
rect -90 282 85 290
rect -64 94 14 124
rect -64 36 -56 94
rect 8 36 14 94
rect -64 28 14 36
rect 43 33 85 282
rect 670 290 9100 332
rect 9141 319 9171 543
rect 670 288 1928 290
rect 670 128 718 288
rect 652 126 730 128
rect 650 118 736 126
rect 124 102 208 112
rect 124 44 138 102
rect 194 78 208 102
rect 194 46 594 78
rect 194 44 208 46
rect -300 -308 -174 -278
rect -300 -372 -274 -308
rect -206 -372 -174 -308
rect -300 -400 -174 -372
rect 47 -465 81 33
rect 124 32 208 44
rect 566 -68 594 46
rect 650 48 656 118
rect 730 48 736 118
rect 1020 110 1078 126
rect 1014 106 1084 110
rect 1014 54 1022 106
rect 1074 94 1084 106
rect 1074 56 1468 94
rect 2512 76 2550 290
rect 3112 104 3198 124
rect 1074 54 1388 56
rect 1014 48 1388 54
rect 650 40 736 48
rect 1374 -10 1388 48
rect 1458 -10 1468 56
rect 1374 -20 1468 -10
rect 2480 46 2592 76
rect 2480 -32 2498 46
rect 2586 -32 2592 46
rect 3112 48 3128 104
rect 3186 48 3198 104
rect 4636 62 4674 290
rect 5222 110 5314 126
rect 3112 36 3198 48
rect 4586 36 4704 62
rect 5222 52 5238 110
rect 5298 52 5314 110
rect 6752 52 6794 290
rect 7338 112 7432 128
rect 7338 56 7352 112
rect 7416 56 7432 112
rect 8882 60 8924 290
rect 9141 289 9511 319
rect 9481 122 9511 289
rect 9454 110 9536 122
rect 5222 44 5314 52
rect 1096 -52 1182 -42
rect 2480 -46 2592 -32
rect 3204 -46 3290 -38
rect 1096 -68 1102 -52
rect 566 -102 1102 -68
rect -722 -680 -618 -662
rect -722 -734 -702 -680
rect -630 -734 -618 -680
rect -722 -752 -618 -734
rect -698 -1182 -662 -752
rect 49 -868 80 -465
rect 566 -625 600 -102
rect 1096 -114 1102 -102
rect 1164 -114 1182 -52
rect 1096 -122 1182 -114
rect 3204 -114 3210 -46
rect 3278 -114 3290 -46
rect 4586 -44 4608 36
rect 4686 -44 4704 36
rect 6724 36 6814 52
rect 7338 42 7432 56
rect 6724 -34 6738 36
rect 6804 -34 6814 36
rect 8840 38 8946 60
rect 4586 -58 4704 -44
rect 5306 -46 5398 -34
rect 3204 -120 3290 -114
rect 5306 -116 5316 -46
rect 5394 -116 5398 -46
rect 6724 -52 6814 -34
rect 7414 -36 7520 -24
rect 648 -144 740 -138
rect 648 -222 662 -144
rect 736 -222 740 -144
rect 648 -230 740 -222
rect 1126 -150 1164 -122
rect 680 -428 730 -230
rect 1126 -262 1162 -150
rect 3232 -262 3268 -120
rect 5306 -122 5398 -116
rect 7414 -112 7430 -36
rect 7502 -112 7520 -36
rect 8840 -36 8860 38
rect 8932 -36 8946 38
rect 9454 46 9466 110
rect 9524 46 9536 110
rect 9454 36 9536 46
rect 8840 -50 8946 -36
rect 7414 -122 7520 -112
rect 1126 -264 3268 -262
rect 5354 -264 5390 -122
rect 1126 -266 5390 -264
rect 7458 -266 7494 -122
rect 1126 -298 9510 -266
rect 680 -466 1760 -428
rect 1282 -504 1392 -494
rect 1282 -572 1302 -504
rect 1384 -572 1392 -504
rect 1282 -586 1392 -572
rect 1012 -620 1090 -606
rect 1012 -625 1024 -620
rect 566 -659 1024 -625
rect 1012 -672 1024 -659
rect 1076 -672 1090 -620
rect 1012 -680 1090 -672
rect 1724 -626 1760 -466
rect 3148 -602 3184 -298
rect 3232 -300 9510 -298
rect 3502 -452 3618 -432
rect 3502 -514 3516 -452
rect 3600 -514 3618 -452
rect 3502 -526 3618 -514
rect 5272 -588 5308 -300
rect 5354 -302 9510 -300
rect 5630 -444 5734 -424
rect 5630 -508 5646 -444
rect 5720 -508 5734 -444
rect 5630 -530 5734 -508
rect 7388 -584 7424 -302
rect 7456 -454 7566 -424
rect 7456 -514 7480 -454
rect 7548 -492 7566 -454
rect 7548 -514 8288 -492
rect 7456 -530 8288 -514
rect 3128 -618 3214 -602
rect 1724 -652 1812 -626
rect 222 -698 344 -686
rect 222 -760 238 -698
rect 338 -760 344 -698
rect 222 -766 344 -760
rect 710 -704 828 -692
rect 222 -770 532 -766
rect 264 -812 532 -770
rect 710 -780 726 -704
rect 810 -780 828 -704
rect 710 -800 828 -780
rect 1122 -726 1234 -708
rect 1122 -786 1138 -726
rect 1208 -786 1234 -726
rect 1724 -710 1746 -652
rect 1808 -710 1812 -652
rect 3128 -670 3146 -618
rect 3198 -670 3214 -618
rect 5246 -608 5330 -588
rect 3128 -684 3214 -670
rect 3844 -644 3934 -624
rect 1724 -728 1812 -710
rect 2832 -702 2948 -688
rect 1122 -802 1234 -786
rect 49 -899 387 -868
rect -306 -992 -178 -970
rect -306 -1072 -286 -992
rect -198 -1072 -178 -992
rect -306 -1090 -178 -1072
rect -698 -1216 -118 -1182
rect -154 -1374 -118 -1216
rect -14 -1332 82 -1310
rect -14 -1358 4 -1332
rect -256 -1400 -110 -1374
rect -256 -1492 -226 -1400
rect -130 -1492 -110 -1400
rect -256 -1516 -110 -1492
rect -72 -1390 4 -1358
rect 66 -1390 82 -1332
rect -72 -1584 -42 -1390
rect -14 -1406 82 -1390
rect 357 -1379 386 -899
rect 482 -1058 530 -812
rect 1754 -886 1796 -728
rect 2832 -764 2842 -702
rect 2928 -764 2948 -702
rect 2832 -780 2948 -764
rect 3250 -718 3356 -698
rect 3250 -780 3272 -718
rect 3336 -780 3356 -718
rect 3844 -716 3856 -644
rect 3924 -716 3934 -644
rect 5246 -660 5266 -608
rect 5320 -660 5330 -608
rect 7358 -608 7454 -584
rect 5246 -676 5330 -660
rect 5960 -650 6044 -622
rect 3844 -726 3934 -716
rect 4930 -696 5060 -686
rect 3250 -800 3356 -780
rect 1754 -1058 1798 -886
rect 2886 -1058 2920 -1056
rect 3848 -1058 3886 -726
rect 4930 -762 4946 -696
rect 5046 -762 5060 -696
rect 4930 -784 5060 -762
rect 5358 -698 5488 -676
rect 5358 -768 5390 -698
rect 5464 -768 5488 -698
rect 5960 -706 5970 -650
rect 5358 -790 5488 -768
rect 5958 -716 5970 -706
rect 6038 -716 6044 -650
rect 7358 -676 7372 -608
rect 7438 -676 7454 -608
rect 7358 -684 7454 -676
rect 8074 -644 8160 -628
rect 5958 -726 6044 -716
rect 8074 -714 8084 -644
rect 8152 -714 8160 -644
rect 8074 -724 8160 -714
rect 5958 -1058 6002 -726
rect 8102 -1058 8140 -724
rect 8248 -790 8288 -530
rect 9474 -552 9510 -302
rect 9564 -482 9596 676
rect 9564 -516 9685 -482
rect 9474 -578 9608 -552
rect 9474 -678 9490 -578
rect 9586 -678 9608 -578
rect 9474 -690 9608 -678
rect 9651 -755 9685 -516
rect 8248 -824 8794 -790
rect 482 -1096 8140 -1058
rect 8754 -1080 8792 -824
rect 482 -1174 530 -1096
rect 434 -1184 530 -1174
rect 434 -1254 442 -1184
rect 520 -1186 530 -1184
rect 792 -1142 902 -1126
rect 520 -1254 528 -1186
rect 792 -1200 810 -1142
rect 884 -1200 902 -1142
rect 2294 -1172 2400 -1150
rect 792 -1210 902 -1200
rect 1954 -1200 2030 -1194
rect 434 -1268 528 -1254
rect 1954 -1266 1962 -1200
rect 2028 -1266 2030 -1200
rect 1954 -1298 2030 -1266
rect 2294 -1246 2310 -1172
rect 2386 -1246 2400 -1172
rect 2886 -1184 2920 -1096
rect 2294 -1268 2400 -1246
rect 2828 -1186 2920 -1184
rect 2828 -1246 2836 -1186
rect 2906 -1246 2920 -1186
rect 3228 -1136 3320 -1124
rect 3228 -1194 3244 -1136
rect 3306 -1194 3320 -1136
rect 4674 -1172 4774 -1154
rect 3228 -1208 3320 -1194
rect 2828 -1252 2920 -1246
rect 4344 -1214 4424 -1194
rect 2000 -1362 2030 -1298
rect 4344 -1282 4356 -1214
rect 4422 -1282 4424 -1214
rect 4674 -1240 4690 -1172
rect 4760 -1240 4774 -1172
rect 5220 -1178 5254 -1096
rect 5864 -1098 6022 -1096
rect 7622 -1098 8140 -1096
rect 5576 -1136 5682 -1126
rect 4674 -1256 4774 -1240
rect 5218 -1182 5314 -1178
rect 5218 -1248 5226 -1182
rect 5294 -1248 5314 -1182
rect 5576 -1200 5594 -1136
rect 5672 -1200 5682 -1136
rect 7076 -1170 7198 -1150
rect 7624 -1166 7658 -1098
rect 8730 -1106 8832 -1080
rect 8730 -1162 8748 -1106
rect 8806 -1162 8832 -1106
rect 5576 -1210 5682 -1200
rect 6734 -1208 6816 -1196
rect 5218 -1254 5314 -1248
rect 4344 -1300 4424 -1282
rect 6734 -1276 6738 -1208
rect 6812 -1276 6816 -1208
rect 7076 -1256 7094 -1170
rect 7184 -1256 7198 -1170
rect 7076 -1274 7198 -1256
rect 7616 -1184 7700 -1166
rect 8730 -1172 8832 -1162
rect 7616 -1254 7622 -1184
rect 7694 -1254 7700 -1184
rect 7616 -1260 7700 -1254
rect 9130 -1202 9204 -1192
rect 9130 -1264 9136 -1202
rect 9198 -1264 9204 -1202
rect 1971 -1368 2030 -1362
rect 2328 -1336 2524 -1308
rect 2328 -1368 2356 -1336
rect 1971 -1379 2356 -1368
rect 357 -1400 2356 -1379
rect 2388 -1384 2466 -1366
rect 357 -1408 2000 -1400
rect 2388 -1436 2398 -1384
rect 2452 -1436 2466 -1384
rect 2496 -1368 2524 -1336
rect 4392 -1368 4424 -1300
rect 4714 -1316 4928 -1288
rect 6734 -1300 6816 -1276
rect 4714 -1368 4742 -1316
rect 2496 -1400 4742 -1368
rect 4778 -1352 4862 -1344
rect 4778 -1418 4784 -1352
rect 4854 -1418 4862 -1352
rect 4900 -1368 4928 -1316
rect 6784 -1368 6816 -1300
rect 9130 -1296 9204 -1264
rect 7110 -1342 7310 -1310
rect 7110 -1368 7144 -1342
rect 4900 -1400 7144 -1368
rect 7272 -1368 7310 -1342
rect 9130 -1368 9160 -1296
rect 4778 -1426 4862 -1418
rect 2388 -1462 2466 -1436
rect 2406 -1490 2450 -1462
rect 4794 -1490 4840 -1426
rect 7172 -1466 7244 -1380
rect 7272 -1400 9160 -1368
rect 2406 -1530 4586 -1490
rect -72 -1612 4390 -1584
rect 4362 -1620 4390 -1612
rect 4546 -1606 4586 -1530
rect 4794 -1536 7146 -1490
rect 7196 -1494 7228 -1466
rect 9652 -1494 9684 -755
rect 7196 -1526 9684 -1494
rect 4362 -1634 4466 -1620
rect 4362 -1648 4394 -1634
rect 4384 -1692 4394 -1648
rect 4458 -1692 4466 -1634
rect 4546 -1636 4736 -1606
rect 4546 -1646 4628 -1636
rect 4384 -1704 4466 -1692
rect 4596 -1704 4628 -1646
rect 4708 -1704 4736 -1636
rect 4596 -1740 4736 -1704
rect 6918 -1620 7036 -1604
rect 7106 -1612 7144 -1536
rect 6918 -1692 6932 -1620
rect 7020 -1692 7036 -1620
rect 6918 -1706 7036 -1692
rect 7074 -1628 7176 -1612
rect 7074 -1682 7100 -1628
rect 7154 -1682 7176 -1628
rect 7074 -1700 7176 -1682
<< via2 >>
rect -536 666 -438 768
rect 7088 664 7158 674
rect 7088 618 7158 664
rect 1500 438 1558 448
rect 1500 392 1502 438
rect 1502 392 1554 438
rect 1554 392 1558 438
rect 2396 428 2462 484
rect 3886 426 3944 432
rect 3886 374 3940 426
rect 3940 374 3944 426
rect 6278 372 6342 428
rect -56 92 8 94
rect -56 38 8 92
rect 138 44 194 102
rect -274 -372 -206 -308
rect 3128 102 3186 104
rect 3128 50 3186 102
rect 3128 48 3186 50
rect 5238 52 5292 110
rect 5292 52 5298 110
rect 7352 56 7416 112
rect 1302 -572 1384 -504
rect 3516 -514 3600 -452
rect 5646 -508 5720 -444
rect 726 -780 810 -704
rect 1138 -786 1208 -726
rect -284 -1072 -200 -992
rect -200 -1072 -198 -992
rect -226 -1492 -130 -1400
rect 2842 -764 2928 -702
rect 3272 -780 3336 -718
rect 4946 -762 5046 -696
rect 5390 -768 5464 -698
rect 810 -1200 884 -1142
rect 2310 -1246 2386 -1172
rect 3244 -1194 3306 -1136
rect 4690 -1240 4760 -1172
rect 5594 -1142 5672 -1136
rect 5594 -1200 5664 -1142
rect 5664 -1200 5672 -1142
rect 7094 -1178 7184 -1170
rect 7094 -1252 7098 -1178
rect 7098 -1252 7174 -1178
rect 7174 -1252 7184 -1178
rect 7094 -1256 7184 -1252
rect 4394 -1692 4458 -1634
rect 6932 -1630 7020 -1620
rect 6932 -1682 6946 -1630
rect 6946 -1682 7008 -1630
rect 7008 -1682 7020 -1630
rect 6932 -1692 7020 -1682
<< metal3 >>
rect -566 768 -418 798
rect -566 666 -536 768
rect -438 666 -418 768
rect 4242 714 4922 786
rect 4242 676 4314 714
rect -566 650 -418 666
rect -568 642 -418 650
rect -568 419 -470 642
rect 2400 604 4314 676
rect 4850 676 4922 714
rect 7066 676 7174 686
rect 4850 674 7174 676
rect 4850 618 7088 674
rect 7158 618 7174 674
rect 4850 604 7174 618
rect 2400 524 2460 604
rect 7066 586 7174 604
rect 2368 484 2484 524
rect 1466 448 1584 472
rect -568 321 -199 419
rect 1466 392 1500 448
rect 1558 392 1584 448
rect 2368 428 2396 484
rect 2462 428 2484 484
rect 6262 458 6368 460
rect 2368 416 2484 428
rect 3862 432 3968 454
rect 1466 348 1584 392
rect 3862 374 3886 432
rect 3944 374 3968 432
rect 3862 360 3968 374
rect 6262 428 6370 458
rect 6262 372 6278 428
rect 6342 372 6370 428
rect 6262 364 6370 372
rect 1466 346 3184 348
rect -295 -308 -200 321
rect 1496 288 3184 346
rect -72 112 30 130
rect 100 112 220 128
rect 3122 124 3184 288
rect 3886 344 3968 360
rect 6310 350 6370 364
rect 7374 350 7436 352
rect 3886 284 5300 344
rect 6310 292 7444 350
rect 6312 288 7444 292
rect 5240 130 5300 284
rect 7374 134 7436 288
rect -72 102 220 112
rect -72 94 138 102
rect -72 38 -56 94
rect 8 52 138 94
rect 8 38 30 52
rect -72 18 30 38
rect 100 44 138 52
rect 194 44 220 102
rect 100 20 220 44
rect 3114 104 3198 124
rect 3114 48 3128 104
rect 3186 48 3198 104
rect 3114 36 3198 48
rect 5212 110 5320 130
rect 5212 52 5238 110
rect 5298 52 5320 110
rect 5212 40 5320 52
rect 7330 112 7436 134
rect 7330 56 7352 112
rect 7416 56 7436 112
rect 7330 40 7436 56
rect -295 -372 -274 -308
rect -206 -372 -200 -308
rect -295 -970 -200 -372
rect 3504 -413 3622 -412
rect 2877 -452 3622 -413
rect 5630 -444 5734 -424
rect 2877 -483 3516 -452
rect 1282 -504 1392 -494
rect 1282 -508 1302 -504
rect 826 -572 1302 -508
rect 1384 -572 1392 -504
rect 826 -692 890 -572
rect 1282 -586 1392 -572
rect 2877 -632 2947 -483
rect 3502 -514 3516 -483
rect 3600 -514 3622 -452
rect 3502 -526 3622 -514
rect 4956 -508 5646 -444
rect 5720 -508 5734 -444
rect 4956 -516 5734 -508
rect 2876 -668 2948 -632
rect 710 -704 890 -692
rect 710 -780 726 -704
rect 810 -756 890 -704
rect 2832 -702 2948 -668
rect 4956 -686 5050 -516
rect 5630 -530 5734 -516
rect 4930 -696 5060 -686
rect 1116 -726 1234 -708
rect 810 -780 828 -756
rect 710 -800 828 -780
rect 1116 -786 1138 -726
rect 1208 -786 1234 -726
rect 2832 -764 2842 -702
rect 2928 -764 2948 -702
rect 2832 -780 2948 -764
rect 3250 -718 3356 -698
rect 3250 -780 3272 -718
rect 3336 -780 3356 -718
rect 1116 -802 1234 -786
rect 3250 -800 3356 -780
rect 4930 -762 4946 -696
rect 5046 -762 5060 -696
rect 4930 -784 5060 -762
rect 5358 -698 5488 -676
rect 5358 -768 5390 -698
rect 5464 -768 5488 -698
rect 5358 -790 5488 -768
rect 1116 -860 1184 -802
rect 836 -928 1184 -860
rect -306 -992 -178 -970
rect -306 -1072 -284 -992
rect -198 -1072 -178 -992
rect -306 -1090 -178 -1072
rect 836 -1112 904 -928
rect 3254 -1108 3320 -800
rect 5406 -842 5488 -790
rect 5406 -918 5680 -842
rect 792 -1142 902 -1112
rect 792 -1200 810 -1142
rect 884 -1200 902 -1142
rect 3210 -1136 3322 -1108
rect 792 -1210 902 -1200
rect 2294 -1172 2400 -1150
rect 2294 -1246 2310 -1172
rect 2386 -1246 2400 -1172
rect 3210 -1194 3244 -1136
rect 3306 -1194 3322 -1136
rect 5576 -1136 5680 -918
rect 4674 -1172 4774 -1154
rect 4674 -1186 4690 -1172
rect 3210 -1210 3322 -1194
rect 4478 -1220 4690 -1186
rect -256 -1400 -110 -1374
rect -256 -1492 -226 -1400
rect -130 -1492 -110 -1400
rect -256 -1516 -110 -1492
rect -217 -1582 -111 -1516
rect 2294 -1582 2400 -1246
rect -217 -1688 2400 -1582
rect 4464 -1240 4690 -1220
rect 4760 -1240 4774 -1172
rect 5576 -1200 5594 -1136
rect 5672 -1200 5680 -1136
rect 7076 -1170 7198 -1150
rect 7076 -1172 7094 -1170
rect 5576 -1208 5680 -1200
rect 4464 -1254 4774 -1240
rect 4464 -1620 4544 -1254
rect 4674 -1256 4774 -1254
rect 6920 -1256 7094 -1172
rect 7184 -1256 7198 -1170
rect 6920 -1274 7198 -1256
rect 6920 -1604 7034 -1274
rect 4384 -1634 4544 -1620
rect 4384 -1692 4394 -1634
rect 4458 -1692 4544 -1634
rect 4384 -1704 4544 -1692
rect 6918 -1620 7036 -1604
rect 6918 -1692 6932 -1620
rect 7020 -1692 7036 -1620
rect 6918 -1706 7036 -1692
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697562905
transform 1 0 816 0 -1 206
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_1
timestamp 1697562905
transform 1 0 -472 0 -1 206
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_2
timestamp 1697562905
transform 1 0 -288 0 1 206
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_3
timestamp 1697562905
transform 1 0 448 0 -1 206
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_4
timestamp 1697562905
transform 1 0 172 0 -1 206
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbp_1  sky130_fd_sc_hd__dfbbp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697562905
transform -1 0 4774 0 -1 -976
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  sky130_fd_sc_hd__dfbbp_1_1
timestamp 1697562905
transform 1 0 2380 0 1 206
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  sky130_fd_sc_hd__dfbbp_1_2
timestamp 1697562905
transform 1 0 4772 0 1 206
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  sky130_fd_sc_hd__dfbbp_1_3
timestamp 1697562905
transform 1 0 7164 0 1 206
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  sky130_fd_sc_hd__dfbbp_1_4
timestamp 1697562905
transform 1 0 -12 0 1 206
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  sky130_fd_sc_hd__dfbbp_1_5
timestamp 1697562905
transform -1 0 2382 0 -1 -976
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  sky130_fd_sc_hd__dfbbp_1_6
timestamp 1697562905
transform -1 0 7166 0 -1 -976
box -38 -48 2430 592
use sky130_fd_sc_hd__dfbbp_1  sky130_fd_sc_hd__dfbbp_1_7
timestamp 1697562905
transform -1 0 9558 0 -1 -976
box -38 -48 2430 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697562905
transform 1 0 1092 0 -1 206
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_1
timestamp 1697562905
transform 1 0 5324 0 -1 206
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_2
timestamp 1697562905
transform 1 0 3208 0 -1 206
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_3
timestamp 1697562905
transform 1 0 7440 0 -1 206
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_4
timestamp 1697562905
transform -1 0 9556 0 1 -882
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_6
timestamp 1697562905
transform -1 0 5324 0 1 -882
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_7
timestamp 1697562905
transform -1 0 7440 0 1 -882
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_8
timestamp 1697562905
transform -1 0 1092 0 1 -882
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrbp_1  sky130_fd_sc_hd__dfrbp_1_9
timestamp 1697562905
transform -1 0 3208 0 1 -882
box -38 -48 2154 592
use sky130_fd_sc_hd__inv_1  sky130_fd_sc_hd__inv_1_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1697562905
transform 1 0 -196 0 -1 206
box -38 -48 314 592
<< labels >>
flabel viali -238 442 -238 442 0 FreeSans 400 0 0 0 cmp
port 0 nsew
flabel viali 226 -24 226 -24 0 FreeSans 400 0 0 0 rstb
port 3 nsew
flabel viali 864 -26 864 -26 0 FreeSans 400 0 0 0 start
port 4 nsew
flabel metal1 -246 750 -246 750 0 FreeSans 400 0 0 0 VDD
port 5 nsew
flabel metal1 -428 202 -428 202 0 FreeSans 400 0 0 0 VSS
port 6 nsew
flabel viali 7114 636 7114 636 0 FreeSans 400 0 0 0 dout5
port 13 nsew
flabel viali 9512 632 9512 632 0 FreeSans 400 0 0 0 dout4
port 14 nsew
flabel viali 4726 638 4726 638 0 FreeSans 400 0 0 0 dout6
port 10 nsew
flabel viali 2046 642 2046 642 0 FreeSans 400 0 0 0 doutb7
port 30 nsew
flabel viali 2432 -1416 2432 -1416 0 FreeSans 400 0 0 0 dout1
port 21 nsew
flabel viali 7212 -1414 7212 -1408 0 FreeSans 400 0 0 0 dout3
port 23 nsew
flabel via1 4816 -1386 4816 -1386 0 FreeSans 400 0 0 0 dout2
port 28 nsew
flabel metal1 34 -1422 34 -1422 0 FreeSans 400 0 0 0 dout0
port 20 nsew
flabel space -20 -1286 -20 -1286 0 FreeSans 240 0 0 0 VSUBS
port 35 nsew
flabel viali 9230 568 9230 568 0 FreeSans 400 0 0 0 doutb4
port 36 nsew
flabel via2 1330 -536 1330 -536 0 FreeSans 400 0 0 0 q5
flabel via2 1186 -760 1186 -760 0 FreeSans 400 0 0 0 nq5
flabel via1 1784 -678 1784 -678 0 FreeSans 400 0 0 0 rst5
flabel via2 2896 -738 2896 -738 0 FreeSans 400 0 0 0 d5
flabel via1 3154 -646 3154 -646 0 FreeSans 400 0 0 0 clk5
flabel viali -416 -34 -416 -34 0 FreeSans 400 0 0 0 clk
port 2 nsew
flabel viali 2332 644 2332 644 0 FreeSans 400 0 0 0 dout7
port 29 nsew
flabel viali 6940 586 6940 586 0 FreeSans 400 0 0 0 doutb5
port 38 nsew
flabel viali 7496 -1338 7496 -1338 0 FreeSans 400 0 0 0 doutb3
port 26 nsew
flabel viali 5104 -1346 5104 -1346 0 FreeSans 400 0 0 0 doutb2
port 27 nsew
flabel viali 2704 -1352 2704 -1352 0 FreeSans 400 0 0 0 doutb1
port 22 nsew
flabel viali 322 -1342 322 -1342 0 FreeSans 400 0 0 0 doutb0
port 19 nsew
flabel viali 4448 640 4448 640 0 FreeSans 400 0 0 0 doutb6
port 39 nsew
flabel via2 1518 412 1518 412 0 FreeSans 240 0 0 0 nq1
flabel via2 3908 400 3908 400 0 FreeSans 240 0 0 0 nq2
flabel via2 6306 392 6306 392 0 FreeSans 240 0 0 0 nq3
flabel via1 8692 400 8692 400 0 FreeSans 240 0 0 0 nq4
flabel via2 160 70 160 70 0 FreeSans 240 0 0 0 clk_t
flabel viali 7092 -28 7092 -28 0 FreeSans 240 0 0 0 q3
flabel viali 9206 -32 9206 -32 0 FreeSans 240 0 0 0 q4
flabel via1 682 82 682 82 0 FreeSans 240 0 0 0 reset
<< end >>

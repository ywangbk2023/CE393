magic
tech sky130A
magscale 1 2
timestamp 1701908128
<< metal3 >>
rect -19716 18812 -13344 18840
rect -19716 12788 -13428 18812
rect -13364 12788 -13344 18812
rect -19716 12760 -13344 12788
rect -13104 18812 -6732 18840
rect -13104 12788 -6816 18812
rect -6752 12788 -6732 18812
rect -13104 12760 -6732 12788
rect -6492 18812 -120 18840
rect -6492 12788 -204 18812
rect -140 12788 -120 18812
rect -6492 12760 -120 12788
rect 120 18812 6492 18840
rect 120 12788 6408 18812
rect 6472 12788 6492 18812
rect 120 12760 6492 12788
rect 6732 18812 13104 18840
rect 6732 12788 13020 18812
rect 13084 12788 13104 18812
rect 6732 12760 13104 12788
rect 13344 18812 19716 18840
rect 13344 12788 19632 18812
rect 19696 12788 19716 18812
rect 13344 12760 19716 12788
rect -19716 12492 -13344 12520
rect -19716 6468 -13428 12492
rect -13364 6468 -13344 12492
rect -19716 6440 -13344 6468
rect -13104 12492 -6732 12520
rect -13104 6468 -6816 12492
rect -6752 6468 -6732 12492
rect -13104 6440 -6732 6468
rect -6492 12492 -120 12520
rect -6492 6468 -204 12492
rect -140 6468 -120 12492
rect -6492 6440 -120 6468
rect 120 12492 6492 12520
rect 120 6468 6408 12492
rect 6472 6468 6492 12492
rect 120 6440 6492 6468
rect 6732 12492 13104 12520
rect 6732 6468 13020 12492
rect 13084 6468 13104 12492
rect 6732 6440 13104 6468
rect 13344 12492 19716 12520
rect 13344 6468 19632 12492
rect 19696 6468 19716 12492
rect 13344 6440 19716 6468
rect -19716 6172 -13344 6200
rect -19716 148 -13428 6172
rect -13364 148 -13344 6172
rect -19716 120 -13344 148
rect -13104 6172 -6732 6200
rect -13104 148 -6816 6172
rect -6752 148 -6732 6172
rect -13104 120 -6732 148
rect -6492 6172 -120 6200
rect -6492 148 -204 6172
rect -140 148 -120 6172
rect -6492 120 -120 148
rect 120 6172 6492 6200
rect 120 148 6408 6172
rect 6472 148 6492 6172
rect 120 120 6492 148
rect 6732 6172 13104 6200
rect 6732 148 13020 6172
rect 13084 148 13104 6172
rect 6732 120 13104 148
rect 13344 6172 19716 6200
rect 13344 148 19632 6172
rect 19696 148 19716 6172
rect 13344 120 19716 148
rect -19716 -148 -13344 -120
rect -19716 -6172 -13428 -148
rect -13364 -6172 -13344 -148
rect -19716 -6200 -13344 -6172
rect -13104 -148 -6732 -120
rect -13104 -6172 -6816 -148
rect -6752 -6172 -6732 -148
rect -13104 -6200 -6732 -6172
rect -6492 -148 -120 -120
rect -6492 -6172 -204 -148
rect -140 -6172 -120 -148
rect -6492 -6200 -120 -6172
rect 120 -148 6492 -120
rect 120 -6172 6408 -148
rect 6472 -6172 6492 -148
rect 120 -6200 6492 -6172
rect 6732 -148 13104 -120
rect 6732 -6172 13020 -148
rect 13084 -6172 13104 -148
rect 6732 -6200 13104 -6172
rect 13344 -148 19716 -120
rect 13344 -6172 19632 -148
rect 19696 -6172 19716 -148
rect 13344 -6200 19716 -6172
rect -19716 -6468 -13344 -6440
rect -19716 -12492 -13428 -6468
rect -13364 -12492 -13344 -6468
rect -19716 -12520 -13344 -12492
rect -13104 -6468 -6732 -6440
rect -13104 -12492 -6816 -6468
rect -6752 -12492 -6732 -6468
rect -13104 -12520 -6732 -12492
rect -6492 -6468 -120 -6440
rect -6492 -12492 -204 -6468
rect -140 -12492 -120 -6468
rect -6492 -12520 -120 -12492
rect 120 -6468 6492 -6440
rect 120 -12492 6408 -6468
rect 6472 -12492 6492 -6468
rect 120 -12520 6492 -12492
rect 6732 -6468 13104 -6440
rect 6732 -12492 13020 -6468
rect 13084 -12492 13104 -6468
rect 6732 -12520 13104 -12492
rect 13344 -6468 19716 -6440
rect 13344 -12492 19632 -6468
rect 19696 -12492 19716 -6468
rect 13344 -12520 19716 -12492
rect -19716 -12788 -13344 -12760
rect -19716 -18812 -13428 -12788
rect -13364 -18812 -13344 -12788
rect -19716 -18840 -13344 -18812
rect -13104 -12788 -6732 -12760
rect -13104 -18812 -6816 -12788
rect -6752 -18812 -6732 -12788
rect -13104 -18840 -6732 -18812
rect -6492 -12788 -120 -12760
rect -6492 -18812 -204 -12788
rect -140 -18812 -120 -12788
rect -6492 -18840 -120 -18812
rect 120 -12788 6492 -12760
rect 120 -18812 6408 -12788
rect 6472 -18812 6492 -12788
rect 120 -18840 6492 -18812
rect 6732 -12788 13104 -12760
rect 6732 -18812 13020 -12788
rect 13084 -18812 13104 -12788
rect 6732 -18840 13104 -18812
rect 13344 -12788 19716 -12760
rect 13344 -18812 19632 -12788
rect 19696 -18812 19716 -12788
rect 13344 -18840 19716 -18812
<< via3 >>
rect -13428 12788 -13364 18812
rect -6816 12788 -6752 18812
rect -204 12788 -140 18812
rect 6408 12788 6472 18812
rect 13020 12788 13084 18812
rect 19632 12788 19696 18812
rect -13428 6468 -13364 12492
rect -6816 6468 -6752 12492
rect -204 6468 -140 12492
rect 6408 6468 6472 12492
rect 13020 6468 13084 12492
rect 19632 6468 19696 12492
rect -13428 148 -13364 6172
rect -6816 148 -6752 6172
rect -204 148 -140 6172
rect 6408 148 6472 6172
rect 13020 148 13084 6172
rect 19632 148 19696 6172
rect -13428 -6172 -13364 -148
rect -6816 -6172 -6752 -148
rect -204 -6172 -140 -148
rect 6408 -6172 6472 -148
rect 13020 -6172 13084 -148
rect 19632 -6172 19696 -148
rect -13428 -12492 -13364 -6468
rect -6816 -12492 -6752 -6468
rect -204 -12492 -140 -6468
rect 6408 -12492 6472 -6468
rect 13020 -12492 13084 -6468
rect 19632 -12492 19696 -6468
rect -13428 -18812 -13364 -12788
rect -6816 -18812 -6752 -12788
rect -204 -18812 -140 -12788
rect 6408 -18812 6472 -12788
rect 13020 -18812 13084 -12788
rect 19632 -18812 19696 -12788
<< mimcap >>
rect -19676 18760 -13676 18800
rect -19676 12840 -19636 18760
rect -13716 12840 -13676 18760
rect -19676 12800 -13676 12840
rect -13064 18760 -7064 18800
rect -13064 12840 -13024 18760
rect -7104 12840 -7064 18760
rect -13064 12800 -7064 12840
rect -6452 18760 -452 18800
rect -6452 12840 -6412 18760
rect -492 12840 -452 18760
rect -6452 12800 -452 12840
rect 160 18760 6160 18800
rect 160 12840 200 18760
rect 6120 12840 6160 18760
rect 160 12800 6160 12840
rect 6772 18760 12772 18800
rect 6772 12840 6812 18760
rect 12732 12840 12772 18760
rect 6772 12800 12772 12840
rect 13384 18760 19384 18800
rect 13384 12840 13424 18760
rect 19344 12840 19384 18760
rect 13384 12800 19384 12840
rect -19676 12440 -13676 12480
rect -19676 6520 -19636 12440
rect -13716 6520 -13676 12440
rect -19676 6480 -13676 6520
rect -13064 12440 -7064 12480
rect -13064 6520 -13024 12440
rect -7104 6520 -7064 12440
rect -13064 6480 -7064 6520
rect -6452 12440 -452 12480
rect -6452 6520 -6412 12440
rect -492 6520 -452 12440
rect -6452 6480 -452 6520
rect 160 12440 6160 12480
rect 160 6520 200 12440
rect 6120 6520 6160 12440
rect 160 6480 6160 6520
rect 6772 12440 12772 12480
rect 6772 6520 6812 12440
rect 12732 6520 12772 12440
rect 6772 6480 12772 6520
rect 13384 12440 19384 12480
rect 13384 6520 13424 12440
rect 19344 6520 19384 12440
rect 13384 6480 19384 6520
rect -19676 6120 -13676 6160
rect -19676 200 -19636 6120
rect -13716 200 -13676 6120
rect -19676 160 -13676 200
rect -13064 6120 -7064 6160
rect -13064 200 -13024 6120
rect -7104 200 -7064 6120
rect -13064 160 -7064 200
rect -6452 6120 -452 6160
rect -6452 200 -6412 6120
rect -492 200 -452 6120
rect -6452 160 -452 200
rect 160 6120 6160 6160
rect 160 200 200 6120
rect 6120 200 6160 6120
rect 160 160 6160 200
rect 6772 6120 12772 6160
rect 6772 200 6812 6120
rect 12732 200 12772 6120
rect 6772 160 12772 200
rect 13384 6120 19384 6160
rect 13384 200 13424 6120
rect 19344 200 19384 6120
rect 13384 160 19384 200
rect -19676 -200 -13676 -160
rect -19676 -6120 -19636 -200
rect -13716 -6120 -13676 -200
rect -19676 -6160 -13676 -6120
rect -13064 -200 -7064 -160
rect -13064 -6120 -13024 -200
rect -7104 -6120 -7064 -200
rect -13064 -6160 -7064 -6120
rect -6452 -200 -452 -160
rect -6452 -6120 -6412 -200
rect -492 -6120 -452 -200
rect -6452 -6160 -452 -6120
rect 160 -200 6160 -160
rect 160 -6120 200 -200
rect 6120 -6120 6160 -200
rect 160 -6160 6160 -6120
rect 6772 -200 12772 -160
rect 6772 -6120 6812 -200
rect 12732 -6120 12772 -200
rect 6772 -6160 12772 -6120
rect 13384 -200 19384 -160
rect 13384 -6120 13424 -200
rect 19344 -6120 19384 -200
rect 13384 -6160 19384 -6120
rect -19676 -6520 -13676 -6480
rect -19676 -12440 -19636 -6520
rect -13716 -12440 -13676 -6520
rect -19676 -12480 -13676 -12440
rect -13064 -6520 -7064 -6480
rect -13064 -12440 -13024 -6520
rect -7104 -12440 -7064 -6520
rect -13064 -12480 -7064 -12440
rect -6452 -6520 -452 -6480
rect -6452 -12440 -6412 -6520
rect -492 -12440 -452 -6520
rect -6452 -12480 -452 -12440
rect 160 -6520 6160 -6480
rect 160 -12440 200 -6520
rect 6120 -12440 6160 -6520
rect 160 -12480 6160 -12440
rect 6772 -6520 12772 -6480
rect 6772 -12440 6812 -6520
rect 12732 -12440 12772 -6520
rect 6772 -12480 12772 -12440
rect 13384 -6520 19384 -6480
rect 13384 -12440 13424 -6520
rect 19344 -12440 19384 -6520
rect 13384 -12480 19384 -12440
rect -19676 -12840 -13676 -12800
rect -19676 -18760 -19636 -12840
rect -13716 -18760 -13676 -12840
rect -19676 -18800 -13676 -18760
rect -13064 -12840 -7064 -12800
rect -13064 -18760 -13024 -12840
rect -7104 -18760 -7064 -12840
rect -13064 -18800 -7064 -18760
rect -6452 -12840 -452 -12800
rect -6452 -18760 -6412 -12840
rect -492 -18760 -452 -12840
rect -6452 -18800 -452 -18760
rect 160 -12840 6160 -12800
rect 160 -18760 200 -12840
rect 6120 -18760 6160 -12840
rect 160 -18800 6160 -18760
rect 6772 -12840 12772 -12800
rect 6772 -18760 6812 -12840
rect 12732 -18760 12772 -12840
rect 6772 -18800 12772 -18760
rect 13384 -12840 19384 -12800
rect 13384 -18760 13424 -12840
rect 19344 -18760 19384 -12840
rect 13384 -18800 19384 -18760
<< mimcapcontact >>
rect -19636 12840 -13716 18760
rect -13024 12840 -7104 18760
rect -6412 12840 -492 18760
rect 200 12840 6120 18760
rect 6812 12840 12732 18760
rect 13424 12840 19344 18760
rect -19636 6520 -13716 12440
rect -13024 6520 -7104 12440
rect -6412 6520 -492 12440
rect 200 6520 6120 12440
rect 6812 6520 12732 12440
rect 13424 6520 19344 12440
rect -19636 200 -13716 6120
rect -13024 200 -7104 6120
rect -6412 200 -492 6120
rect 200 200 6120 6120
rect 6812 200 12732 6120
rect 13424 200 19344 6120
rect -19636 -6120 -13716 -200
rect -13024 -6120 -7104 -200
rect -6412 -6120 -492 -200
rect 200 -6120 6120 -200
rect 6812 -6120 12732 -200
rect 13424 -6120 19344 -200
rect -19636 -12440 -13716 -6520
rect -13024 -12440 -7104 -6520
rect -6412 -12440 -492 -6520
rect 200 -12440 6120 -6520
rect 6812 -12440 12732 -6520
rect 13424 -12440 19344 -6520
rect -19636 -18760 -13716 -12840
rect -13024 -18760 -7104 -12840
rect -6412 -18760 -492 -12840
rect 200 -18760 6120 -12840
rect 6812 -18760 12732 -12840
rect 13424 -18760 19344 -12840
<< metal4 >>
rect -16728 18761 -16624 18960
rect -13448 18812 -13344 18960
rect -19637 18760 -13715 18761
rect -19637 12840 -19636 18760
rect -13716 12840 -13715 18760
rect -19637 12839 -13715 12840
rect -16728 12441 -16624 12839
rect -13448 12788 -13428 18812
rect -13364 12788 -13344 18812
rect -10116 18761 -10012 18960
rect -6836 18812 -6732 18960
rect -13025 18760 -7103 18761
rect -13025 12840 -13024 18760
rect -7104 12840 -7103 18760
rect -13025 12839 -7103 12840
rect -13448 12492 -13344 12788
rect -19637 12440 -13715 12441
rect -19637 6520 -19636 12440
rect -13716 6520 -13715 12440
rect -19637 6519 -13715 6520
rect -16728 6121 -16624 6519
rect -13448 6468 -13428 12492
rect -13364 6468 -13344 12492
rect -10116 12441 -10012 12839
rect -6836 12788 -6816 18812
rect -6752 12788 -6732 18812
rect -3504 18761 -3400 18960
rect -224 18812 -120 18960
rect -6413 18760 -491 18761
rect -6413 12840 -6412 18760
rect -492 12840 -491 18760
rect -6413 12839 -491 12840
rect -6836 12492 -6732 12788
rect -13025 12440 -7103 12441
rect -13025 6520 -13024 12440
rect -7104 6520 -7103 12440
rect -13025 6519 -7103 6520
rect -13448 6172 -13344 6468
rect -19637 6120 -13715 6121
rect -19637 200 -19636 6120
rect -13716 200 -13715 6120
rect -19637 199 -13715 200
rect -16728 -199 -16624 199
rect -13448 148 -13428 6172
rect -13364 148 -13344 6172
rect -10116 6121 -10012 6519
rect -6836 6468 -6816 12492
rect -6752 6468 -6732 12492
rect -3504 12441 -3400 12839
rect -224 12788 -204 18812
rect -140 12788 -120 18812
rect 3108 18761 3212 18960
rect 6388 18812 6492 18960
rect 199 18760 6121 18761
rect 199 12840 200 18760
rect 6120 12840 6121 18760
rect 199 12839 6121 12840
rect -224 12492 -120 12788
rect -6413 12440 -491 12441
rect -6413 6520 -6412 12440
rect -492 6520 -491 12440
rect -6413 6519 -491 6520
rect -6836 6172 -6732 6468
rect -13025 6120 -7103 6121
rect -13025 200 -13024 6120
rect -7104 200 -7103 6120
rect -13025 199 -7103 200
rect -13448 -148 -13344 148
rect -19637 -200 -13715 -199
rect -19637 -6120 -19636 -200
rect -13716 -6120 -13715 -200
rect -19637 -6121 -13715 -6120
rect -16728 -6519 -16624 -6121
rect -13448 -6172 -13428 -148
rect -13364 -6172 -13344 -148
rect -10116 -199 -10012 199
rect -6836 148 -6816 6172
rect -6752 148 -6732 6172
rect -3504 6121 -3400 6519
rect -224 6468 -204 12492
rect -140 6468 -120 12492
rect 3108 12441 3212 12839
rect 6388 12788 6408 18812
rect 6472 12788 6492 18812
rect 9720 18761 9824 18960
rect 13000 18812 13104 18960
rect 6811 18760 12733 18761
rect 6811 12840 6812 18760
rect 12732 12840 12733 18760
rect 6811 12839 12733 12840
rect 6388 12492 6492 12788
rect 199 12440 6121 12441
rect 199 6520 200 12440
rect 6120 6520 6121 12440
rect 199 6519 6121 6520
rect -224 6172 -120 6468
rect -6413 6120 -491 6121
rect -6413 200 -6412 6120
rect -492 200 -491 6120
rect -6413 199 -491 200
rect -6836 -148 -6732 148
rect -13025 -200 -7103 -199
rect -13025 -6120 -13024 -200
rect -7104 -6120 -7103 -200
rect -13025 -6121 -7103 -6120
rect -13448 -6468 -13344 -6172
rect -19637 -6520 -13715 -6519
rect -19637 -12440 -19636 -6520
rect -13716 -12440 -13715 -6520
rect -19637 -12441 -13715 -12440
rect -16728 -12839 -16624 -12441
rect -13448 -12492 -13428 -6468
rect -13364 -12492 -13344 -6468
rect -10116 -6519 -10012 -6121
rect -6836 -6172 -6816 -148
rect -6752 -6172 -6732 -148
rect -3504 -199 -3400 199
rect -224 148 -204 6172
rect -140 148 -120 6172
rect 3108 6121 3212 6519
rect 6388 6468 6408 12492
rect 6472 6468 6492 12492
rect 9720 12441 9824 12839
rect 13000 12788 13020 18812
rect 13084 12788 13104 18812
rect 16332 18761 16436 18960
rect 19612 18812 19716 18960
rect 13423 18760 19345 18761
rect 13423 12840 13424 18760
rect 19344 12840 19345 18760
rect 13423 12839 19345 12840
rect 13000 12492 13104 12788
rect 6811 12440 12733 12441
rect 6811 6520 6812 12440
rect 12732 6520 12733 12440
rect 6811 6519 12733 6520
rect 6388 6172 6492 6468
rect 199 6120 6121 6121
rect 199 200 200 6120
rect 6120 200 6121 6120
rect 199 199 6121 200
rect -224 -148 -120 148
rect -6413 -200 -491 -199
rect -6413 -6120 -6412 -200
rect -492 -6120 -491 -200
rect -6413 -6121 -491 -6120
rect -6836 -6468 -6732 -6172
rect -13025 -6520 -7103 -6519
rect -13025 -12440 -13024 -6520
rect -7104 -12440 -7103 -6520
rect -13025 -12441 -7103 -12440
rect -13448 -12788 -13344 -12492
rect -19637 -12840 -13715 -12839
rect -19637 -18760 -19636 -12840
rect -13716 -18760 -13715 -12840
rect -19637 -18761 -13715 -18760
rect -16728 -18960 -16624 -18761
rect -13448 -18812 -13428 -12788
rect -13364 -18812 -13344 -12788
rect -10116 -12839 -10012 -12441
rect -6836 -12492 -6816 -6468
rect -6752 -12492 -6732 -6468
rect -3504 -6519 -3400 -6121
rect -224 -6172 -204 -148
rect -140 -6172 -120 -148
rect 3108 -199 3212 199
rect 6388 148 6408 6172
rect 6472 148 6492 6172
rect 9720 6121 9824 6519
rect 13000 6468 13020 12492
rect 13084 6468 13104 12492
rect 16332 12441 16436 12839
rect 19612 12788 19632 18812
rect 19696 12788 19716 18812
rect 19612 12492 19716 12788
rect 13423 12440 19345 12441
rect 13423 6520 13424 12440
rect 19344 6520 19345 12440
rect 13423 6519 19345 6520
rect 13000 6172 13104 6468
rect 6811 6120 12733 6121
rect 6811 200 6812 6120
rect 12732 200 12733 6120
rect 6811 199 12733 200
rect 6388 -148 6492 148
rect 199 -200 6121 -199
rect 199 -6120 200 -200
rect 6120 -6120 6121 -200
rect 199 -6121 6121 -6120
rect -224 -6468 -120 -6172
rect -6413 -6520 -491 -6519
rect -6413 -12440 -6412 -6520
rect -492 -12440 -491 -6520
rect -6413 -12441 -491 -12440
rect -6836 -12788 -6732 -12492
rect -13025 -12840 -7103 -12839
rect -13025 -18760 -13024 -12840
rect -7104 -18760 -7103 -12840
rect -13025 -18761 -7103 -18760
rect -13448 -18960 -13344 -18812
rect -10116 -18960 -10012 -18761
rect -6836 -18812 -6816 -12788
rect -6752 -18812 -6732 -12788
rect -3504 -12839 -3400 -12441
rect -224 -12492 -204 -6468
rect -140 -12492 -120 -6468
rect 3108 -6519 3212 -6121
rect 6388 -6172 6408 -148
rect 6472 -6172 6492 -148
rect 9720 -199 9824 199
rect 13000 148 13020 6172
rect 13084 148 13104 6172
rect 16332 6121 16436 6519
rect 19612 6468 19632 12492
rect 19696 6468 19716 12492
rect 19612 6172 19716 6468
rect 13423 6120 19345 6121
rect 13423 200 13424 6120
rect 19344 200 19345 6120
rect 13423 199 19345 200
rect 13000 -148 13104 148
rect 6811 -200 12733 -199
rect 6811 -6120 6812 -200
rect 12732 -6120 12733 -200
rect 6811 -6121 12733 -6120
rect 6388 -6468 6492 -6172
rect 199 -6520 6121 -6519
rect 199 -12440 200 -6520
rect 6120 -12440 6121 -6520
rect 199 -12441 6121 -12440
rect -224 -12788 -120 -12492
rect -6413 -12840 -491 -12839
rect -6413 -18760 -6412 -12840
rect -492 -18760 -491 -12840
rect -6413 -18761 -491 -18760
rect -6836 -18960 -6732 -18812
rect -3504 -18960 -3400 -18761
rect -224 -18812 -204 -12788
rect -140 -18812 -120 -12788
rect 3108 -12839 3212 -12441
rect 6388 -12492 6408 -6468
rect 6472 -12492 6492 -6468
rect 9720 -6519 9824 -6121
rect 13000 -6172 13020 -148
rect 13084 -6172 13104 -148
rect 16332 -199 16436 199
rect 19612 148 19632 6172
rect 19696 148 19716 6172
rect 19612 -148 19716 148
rect 13423 -200 19345 -199
rect 13423 -6120 13424 -200
rect 19344 -6120 19345 -200
rect 13423 -6121 19345 -6120
rect 13000 -6468 13104 -6172
rect 6811 -6520 12733 -6519
rect 6811 -12440 6812 -6520
rect 12732 -12440 12733 -6520
rect 6811 -12441 12733 -12440
rect 6388 -12788 6492 -12492
rect 199 -12840 6121 -12839
rect 199 -18760 200 -12840
rect 6120 -18760 6121 -12840
rect 199 -18761 6121 -18760
rect -224 -18960 -120 -18812
rect 3108 -18960 3212 -18761
rect 6388 -18812 6408 -12788
rect 6472 -18812 6492 -12788
rect 9720 -12839 9824 -12441
rect 13000 -12492 13020 -6468
rect 13084 -12492 13104 -6468
rect 16332 -6519 16436 -6121
rect 19612 -6172 19632 -148
rect 19696 -6172 19716 -148
rect 19612 -6468 19716 -6172
rect 13423 -6520 19345 -6519
rect 13423 -12440 13424 -6520
rect 19344 -12440 19345 -6520
rect 13423 -12441 19345 -12440
rect 13000 -12788 13104 -12492
rect 6811 -12840 12733 -12839
rect 6811 -18760 6812 -12840
rect 12732 -18760 12733 -12840
rect 6811 -18761 12733 -18760
rect 6388 -18960 6492 -18812
rect 9720 -18960 9824 -18761
rect 13000 -18812 13020 -12788
rect 13084 -18812 13104 -12788
rect 16332 -12839 16436 -12441
rect 19612 -12492 19632 -6468
rect 19696 -12492 19716 -6468
rect 19612 -12788 19716 -12492
rect 13423 -12840 19345 -12839
rect 13423 -18760 13424 -12840
rect 19344 -18760 19345 -12840
rect 13423 -18761 19345 -18760
rect 13000 -18960 13104 -18812
rect 16332 -18960 16436 -18761
rect 19612 -18812 19632 -12788
rect 19696 -18812 19716 -12788
rect 19612 -18960 19716 -18812
<< properties >>
string FIXED_BBOX 13344 12760 19424 18840
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 30 l 30 val 1.822k carea 2.00 cperi 0.19 nx 6 ny 6 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>

* NGSPICE file created from SARLOGIC_top.ext - technology: sky130A

.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.115 pd=1.08 as=0.205 ps=2.1 w=0.79 l=0.15
X1 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.205 pd=2.1 as=0.115 ps=1.08 w=0.79 l=0.15
X3 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.135 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N a_2136_47#
X0 a_788_47# a_942_21# a_648_21# VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 VPWR RESET_B a_942_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X2 VGND a_1429_21# a_1364_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.066 ps=0.745 w=0.42 l=0.15
X3 VPWR a_942_21# a_1663_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.218 pd=2.2 as=0.0882 ps=1.05 w=0.84 l=0.15
X4 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.109 ps=1.36 w=0.42 l=0.15
X6 VPWR a_1429_21# a_1341_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0924 ps=0.86 w=0.42 l=0.15
X7 a_474_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X8 a_1545_47# a_942_21# a_1429_21# VNB sky130_fd_pr__nfet_01v8 ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9 VPWR a_1429_21# a_2136_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.33 as=0.166 ps=1.8 w=0.64 l=0.15
X10 a_582_47# a_193_47# a_474_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0671 pd=0.75 as=0.0684 ps=0.74 w=0.36 l=0.15
X11 a_1429_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.123 pd=1.17 as=0.0819 ps=0.81 w=0.42 l=0.15
X12 a_648_21# a_474_413# a_788_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.101 ps=0.99 w=0.64 l=0.15
X13 a_1341_413# a_193_47# a_1255_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0924 pd=0.86 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 a_1663_329# a_1255_47# a_1429_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=1.05 as=0.123 ps=1.17 w=0.84 l=0.15
X15 a_1160_47# a_648_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.166 ps=1.8 w=0.64 l=0.15
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 a_1255_47# a_27_47# a_1113_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.174 ps=1.41 w=0.42 l=0.15
X18 Q a_2136_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.33 w=1 l=0.15
X19 a_648_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.147 pd=1.23 as=0.0798 ps=0.8 w=0.42 l=0.15
X20 a_788_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.101 pd=0.99 as=0.084 ps=0.82 w=0.42 l=0.15
X21 Q_N a_1429_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X22 VGND RESET_B a_942_21# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X23 Q a_2136_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X24 VPWR a_942_21# a_892_329# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.225 pd=1.38 as=0.113 ps=1.11 w=0.84 l=0.15
X25 a_558_413# a_27_47# a_474_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 VGND a_648_21# a_582_47# VNB sky130_fd_pr__nfet_01v8 ad=0.084 pd=0.82 as=0.0671 ps=0.75 w=0.42 l=0.15
X27 a_892_329# a_474_413# a_648_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.113 pd=1.11 as=0.147 ps=1.23 w=0.84 l=0.15
X28 VGND a_1429_21# a_2136_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.109 ps=1.36 w=0.42 l=0.15
X29 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X30 a_474_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0662 ps=0.735 w=0.42 l=0.15
X31 a_1364_47# a_27_47# a_1255_47# VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0711 ps=0.755 w=0.36 l=0.15
X32 a_1255_47# a_193_47# a_1160_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0935 ps=0.965 w=0.36 l=0.15
X33 Q_N a_1429_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X34 a_1545_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.12 pd=1.08 as=0.0588 ps=0.7 w=0.42 l=0.15
X35 VPWR a_648_21# a_558_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X36 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.109 ps=1.36 w=0.42 l=0.15
X37 a_1113_329# a_648_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.174 pd=1.41 as=0.225 ps=1.38 w=0.84 l=0.15
X38 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X39 a_1429_21# a_1255_47# a_1545_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0864 pd=0.91 as=0.12 ps=1.08 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrbp_1 CLK D RESET_B VGND VNB VPB VPWR Q Q_N a_1847_47#
+ a_27_47#
X0 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.213 ps=1.67 w=1 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.14 ps=1.1 w=0.42 l=0.15
X3 VPWR a_1283_21# a_1847_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.34 as=0.166 ps=1.8 w=0.64 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.064 ps=0.725 w=0.42 l=0.15
X6 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.116 pd=0.97 as=0.0724 ps=0.765 w=0.42 l=0.15
X7 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.135 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X8 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.166 ps=1.8 w=0.64 l=0.15
X9 Q_N a_1847_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1 ps=0.985 w=0.65 l=0.15
X10 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.109 ps=1.36 w=0.42 l=0.15
X11 VGND a_1283_21# a_1847_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1 pd=0.985 as=0.109 ps=1.36 w=0.42 l=0.15
X12 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.135 ps=1.15 w=0.64 l=0.15
X13 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X14 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.109 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X15 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.129 ps=1.18 w=0.42 l=0.15
X16 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X17 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.064 pd=0.725 as=0.125 ps=1.01 w=0.42 l=0.15
X18 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0724 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X19 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.221 ps=1.89 w=0.42 l=0.15
X20 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X21 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.213 pd=1.67 as=0.0567 ps=0.69 w=0.42 l=0.15
X22 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.166 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0703 pd=0.755 as=0.116 ps=0.97 w=0.42 l=0.15
X26 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__nfet_01v8 ad=0.14 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X27 Q_N a_1847_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.34 w=1 l=0.15
X28 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.01 as=0.0669 ps=0.75 w=0.42 l=0.15
X29 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.109 pd=1.36 as=0.0703 ps=0.755 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.109 ps=1.36 w=0.42 l=0.15
X31 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.129 pd=1.18 as=0.218 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_fd_sc_hd__inv_1 A VGND VNB VPB VPWR Y
X0 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
.ends

.subckt SARLOGIC_layout cmp clk rstb start VDD VSS dout6 dout5 dout4 doutb0 dout0
+ dout1 doutb1 dout3 doutb3 doutb2 dout2 dout7 doutb7 doutb4 doutb5 doutb6 VSUBS
Xsky130_fd_sc_hd__buf_1_4 rstb VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB VDD sky130_fd_sc_hd__buf_1_4/X
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__dfbbp_1_0 dout0 sky130_fd_sc_hd__buf_1_2/X rst5 sky130_fd_sc_hd__dfrbp_1_6/Q_N
+ VSS VSUBS sky130_fd_sc_hd__dfbbp_1_7/VPB VDD dout1 doutb1 sky130_fd_sc_hd__dfbbp_1_0/a_2136_47#
+ sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_1 dout5 sky130_fd_sc_hd__buf_1_2/X rst5 nq2 VSS VSUBS sky130_fd_sc_hd__buf_1_2/VPB
+ VDD dout6 doutb6 sky130_fd_sc_hd__dfbbp_1_1/a_2136_47# sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_2 dout4 sky130_fd_sc_hd__buf_1_2/X rst5 nq3 VSS VSUBS sky130_fd_sc_hd__buf_1_2/VPB
+ VDD dout5 sky130_fd_sc_hd__dfbbp_1_2/Q_N doutb5 sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_3 sky130_fd_sc_hd__dfbbp_1_3/CLK sky130_fd_sc_hd__buf_1_2/X
+ rst5 nq4 VSS VSUBS sky130_fd_sc_hd__buf_1_2/VPB VDD dout4 doutb4 sky130_fd_sc_hd__dfbbp_1_3/a_2136_47#
+ sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_4 dout6 sky130_fd_sc_hd__buf_1_2/X rst5 nq1 VSS VSUBS sky130_fd_sc_hd__buf_1_2/VPB
+ VDD dout7 doutb7 sky130_fd_sc_hd__dfbbp_1_4/a_2136_47# sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_6 dout1 sky130_fd_sc_hd__buf_1_2/X rst5 sky130_fd_sc_hd__dfrbp_1_7/Q_N
+ VSS VSUBS sky130_fd_sc_hd__dfbbp_1_7/VPB VDD sky130_fd_sc_hd__dfbbp_1_6/Q doutb2
+ sky130_fd_sc_hd__dfbbp_1_6/a_2136_47# sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_5 sky130_fd_sc_hd__dfrbp_1_8/Q sky130_fd_sc_hd__buf_1_2/X
+ rst5 nq5 VSS VSUBS sky130_fd_sc_hd__dfbbp_1_7/VPB VDD dout0 doutb0 sky130_fd_sc_hd__dfbbp_1_5/a_2136_47#
+ sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfbbp_1_7 dout2 sky130_fd_sc_hd__buf_1_2/X rst5 sky130_fd_sc_hd__dfrbp_1_4/Q_N
+ VSS VSUBS sky130_fd_sc_hd__dfbbp_1_7/VPB VDD dout3 doutb3 sky130_fd_sc_hd__dfbbp_1_7/a_2136_47#
+ sky130_fd_sc_hd__dfbbp_1
Xsky130_fd_sc_hd__dfrbp_1_0 clk5 sky130_fd_sc_hd__buf_1_0/X rst5 VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ VDD sky130_fd_sc_hd__dfrbp_1_2/D nq1 sky130_fd_sc_hd__dfrbp_1_0/a_1847_47# sky130_fd_sc_hd__buf_1_0/X
+ sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_1 clk5 sky130_fd_sc_hd__dfrbp_1_2/Q rst5 VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ VDD q3 nq3 sky130_fd_sc_hd__dfrbp_1_1/a_1847_47# sky130_fd_sc_hd__dfrbp_1_1/a_27_47#
+ sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_2 clk5 sky130_fd_sc_hd__dfrbp_1_2/D rst5 VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ VDD sky130_fd_sc_hd__dfrbp_1_2/Q nq2 sky130_fd_sc_hd__dfrbp_1_2/a_1847_47# sky130_fd_sc_hd__dfrbp_1_2/a_27_47#
+ sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_3 clk5 q3 rst5 VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB VDD
+ q4 nq4 sky130_fd_sc_hd__dfrbp_1_3/a_1847_47# sky130_fd_sc_hd__dfrbp_1_3/a_27_47#
+ sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_4 clk5 q4 rst5 VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB VDD
+ sky130_fd_sc_hd__dfrbp_1_7/D sky130_fd_sc_hd__dfrbp_1_4/Q_N sky130_fd_sc_hd__dfrbp_1_4/a_1847_47#
+ sky130_fd_sc_hd__dfrbp_1_4/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_6 clk5 sky130_fd_sc_hd__dfrbp_1_7/Q rst5 VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ VDD d5 sky130_fd_sc_hd__dfrbp_1_6/Q_N sky130_fd_sc_hd__dfrbp_1_6/a_1847_47# sky130_fd_sc_hd__dfrbp_1_6/a_27_47#
+ sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__dfrbp_1_7 clk5 sky130_fd_sc_hd__dfrbp_1_7/D rst5 VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ VDD sky130_fd_sc_hd__dfrbp_1_7/Q sky130_fd_sc_hd__dfrbp_1_7/Q_N sky130_fd_sc_hd__dfrbp_1_7/a_1847_47#
+ sky130_fd_sc_hd__dfrbp_1_7/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__buf_1_0 start VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB VDD sky130_fd_sc_hd__buf_1_0/X
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__dfrbp_1_8 sky130_fd_sc_hd__dfrbp_1_8/CLK q5 rst5 VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ VDD sky130_fd_sc_hd__dfrbp_1_8/Q sky130_fd_sc_hd__dfrbp_1_8/Q_N sky130_fd_sc_hd__dfrbp_1_8/a_1847_47#
+ sky130_fd_sc_hd__dfrbp_1_8/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__inv_1_0 sky130_fd_sc_hd__inv_1_0/A VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ VDD clk5 sky130_fd_sc_hd__inv_1
Xsky130_fd_sc_hd__buf_1_1 clk VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB VDD sky130_fd_sc_hd__inv_1_0/A
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__dfrbp_1_9 clk5 d5 rst5 VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB VDD
+ sky130_fd_sc_hd__dfrbp_1_9/Q nq5 q5 sky130_fd_sc_hd__dfrbp_1_9/a_27_47# sky130_fd_sc_hd__dfrbp_1
Xsky130_fd_sc_hd__buf_1_2 cmp VSS VSUBS sky130_fd_sc_hd__buf_1_2/VPB VDD sky130_fd_sc_hd__buf_1_2/X
+ sky130_fd_sc_hd__buf_1
Xsky130_fd_sc_hd__buf_1_3 sky130_fd_sc_hd__buf_1_4/X VSS VSUBS sky130_fd_sc_hd__inv_1_0/VPB
+ VDD rst5 sky130_fd_sc_hd__buf_1
.ends

.subckt SARLOGIC_top
XSARLOGIC_layout_0 SARLOGIC_layout_0/cmp SARLOGIC_layout_0/clk SARLOGIC_layout_0/rstb
+ SARLOGIC_layout_0/start SARLOGIC_layout_0/VDD SARLOGIC_layout_0/VSS SARLOGIC_layout_0/dout6
+ SARLOGIC_layout_0/dout5 SARLOGIC_layout_0/dout4 SARLOGIC_layout_0/doutb0 SARLOGIC_layout_0/dout0
+ SARLOGIC_layout_0/dout1 SARLOGIC_layout_0/doutb1 SARLOGIC_layout_0/dout3 SARLOGIC_layout_0/doutb3
+ SARLOGIC_layout_0/doutb2 SARLOGIC_layout_0/dout2 SARLOGIC_layout_0/dout7 SARLOGIC_layout_0/doutb7
+ SARLOGIC_layout_0/doutb4 SARLOGIC_layout_0/doutb5 SARLOGIC_layout_0/doutb6 VSUBS
+ SARLOGIC_layout
.ends

